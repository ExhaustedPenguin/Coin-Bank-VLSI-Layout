* File: Coin_bank.pex.sp
* Created: Sat Jan 20 20:42:00 2024
* Program "Calibre xRC"
* Version "v2021.3_35.19"
* 
.include "Coin_bank.pex.sp.pex"
.subckt COIN_BANK  CLK STATE0 STORE STATE1 INIT3 INIT2 INIT1 POWER INIT0 S1 VSS
+ VDD M3 M1 M2 M0 S0 S3 S2 MO1 MO3 MO0 MO2
* 
* MO2	MO2
* MO0	MO0
* MO3	MO3
* MO1	MO1
* S2	S2
* S3	S3
* S0	S0
* M0	M0
* M2	M2
* M1	M1
* M3	M3
* VDD	VDD
* VSS	VSS
* S1	S1
* INIT0	INIT0
* POWER	POWER
* INIT1	INIT1
* INIT2	INIT2
* INIT3	INIT3
* STATE1	STATE1
* STORE	STORE
* STATE0	STATE0
* CLK	CLK
M0 N_VSS_M0_d N_6_M0_g N_49_M0_s N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06
+ AD=1.395e-12 AS=2.85e-12 PD=9.3e-07 PS=4.9e-06
M1 N_5_M1_d N_49_M1_g N_VSS_M1_s N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06
+ AD=1.395e-12 AS=2.7e-12 PD=9.3e-07 PS=4.8e-06
M2 N_49_M2_d N_50_M2_g N_VSS_M2_s N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06
+ AD=1.395e-12 AS=1.395e-12 PD=9.3e-07 PS=9.3e-07
M3 N_VSS_M3_d N_26_M3_g N_5_M3_s N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06
+ AD=2.82e-12 AS=1.395e-12 PD=4.88e-06 PS=9.3e-07
M4 N_VSS_M4_d N_STATE1_M4_g N_49_M4_s N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06
+ AD=2.82e-12 AS=1.395e-12 PD=4.88e-06 PS=9.3e-07
M5 N_68_M5_d N_STORE_M5_g N_VSS_M5_s N_VSS_X24/M0_b N_18 L=1.8e-07 W=9e-06
+ AD=4.185e-12 AS=8.46e-12 PD=9.3e-07 PS=1.088e-05
M6 N_69_M6_d N_11_M6_g N_68_M6_s N_VSS_X24/M0_b N_18 L=1.8e-07 W=9e-06
+ AD=4.185e-12 AS=4.185e-12 PD=9.3e-07 PS=9.3e-07
M7 N_70_M7_d N_STATE0_M7_g N_69_M7_s N_VSS_X24/M0_b N_18 L=1.8e-07 W=9e-06
+ AD=3.915e-12 AS=4.185e-12 PD=8.7e-07 PS=9.3e-07
M8 N_51_M8_d N_POWER_M8_g N_70_M8_s N_VSS_X24/M0_b N_18 L=1.8e-07 W=9e-06
+ AD=6.66e-12 AS=3.915e-12 PD=1.048e-05 PS=8.7e-07
M9 N_71_M9_d N_POWER_M9_g N_29_M9_s N_VSS_X24/M0_b N_18 L=1.8e-07 W=9e-06
+ AD=4.185e-12 AS=8.55e-12 PD=9.3e-07 PS=1.09e-05
M10 N_72_M10_d N_STATE1_M10_g N_71_M10_s N_VSS_X24/M0_b N_18 L=1.8e-07 W=9e-06
+ AD=4.185e-12 AS=4.185e-12 PD=9.3e-07 PS=9.3e-07
M11 N_VSS_M11_d N_6_M11_g N_72_M11_s N_VSS_X24/M0_b N_18 L=1.8e-07 W=9e-06
+ AD=8.46e-12 AS=4.185e-12 PD=1.088e-05 PS=9.3e-07
M12 N_65_M12_d N_6_M12_g N_49_M12_s N_VDD_M12_b P_18 L=1.8e-07 W=6e-06
+ AD=2.79e-12 AS=5.7e-12 PD=9.3e-07 PS=7.9e-06
M13 N_66_M13_d N_49_M13_g N_5_M13_s N_VDD_M13_b P_18 L=1.8e-07 W=6e-06
+ AD=2.79e-12 AS=5.4e-12 PD=9.3e-07 PS=7.8e-06
M14 N_67_M14_d N_50_M14_g N_65_M14_s N_VDD_M12_b P_18 L=1.8e-07 W=6e-06
+ AD=2.79e-12 AS=2.79e-12 PD=9.3e-07 PS=9.3e-07
M15 N_VDD_M15_d N_26_M15_g N_66_M15_s N_VDD_M13_b P_18 L=1.8e-07 W=6e-06
+ AD=5.64e-12 AS=2.79e-12 PD=7.88e-06 PS=9.3e-07
M16 N_VDD_M16_d N_STATE1_M16_g N_67_M16_s N_VDD_M12_b P_18 L=1.8e-07 W=6e-06
+ AD=5.64e-12 AS=2.79e-12 PD=7.88e-06 PS=9.3e-07
M17 N_VDD_M17_d N_STORE_M17_g N_51_M17_s N_VDD_M17_b P_18 L=1.8e-07 W=6e-06
+ AD=2.79e-12 AS=5.64e-12 PD=9.3e-07 PS=7.88e-06
M18 N_51_M18_d N_11_M18_g N_VDD_M18_s N_VDD_M17_b P_18 L=1.8e-07 W=6e-06
+ AD=2.79e-12 AS=2.79e-12 PD=9.3e-07 PS=9.3e-07
M19 N_VDD_M19_d N_STATE0_M19_g N_51_M19_s N_VDD_M17_b P_18 L=1.8e-07 W=6e-06
+ AD=2.61e-12 AS=2.79e-12 PD=8.7e-07 PS=9.3e-07
M20 N_51_M20_d N_POWER_M20_g N_VDD_M20_s N_VDD_M17_b P_18 L=1.8e-07 W=6e-06
+ AD=4.44e-12 AS=2.61e-12 PD=7.48e-06 PS=8.7e-07
M21 N_VDD_M21_d N_POWER_M21_g N_29_M21_s N_VDD_M21_b P_18 L=1.8e-07 W=6e-06
+ AD=2.79e-12 AS=5.7e-12 PD=9.3e-07 PS=7.9e-06
M22 N_29_M22_d N_STATE1_M22_g N_VDD_M22_s N_VDD_M21_b P_18 L=1.8e-07 W=6e-06
+ AD=2.79e-12 AS=2.79e-12 PD=9.3e-07 PS=9.3e-07
M23 N_VDD_M23_d N_6_M23_g N_29_M23_s N_VDD_M21_b P_18 L=1.8e-07 W=6e-06
+ AD=5.64e-12 AS=2.79e-12 PD=7.88e-06 PS=9.3e-07
mX24/M0 N_X24/6_X24/M0_d N_34_X24/M0_g N_VSS_X24/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07 PS=7.88e-06
mX24/M1 N_27_X24/M1_d N_28_X24/M1_g N_X24/6_X24/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06 PS=9.3e-07
mX24/M2 N_27_X24/M2_d N_34_X24/M2_g N_VDD_X24/M2_s N_VDD_X24/M2_b P_18 L=1.8e-07
+ W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07 PS=7.88e-06
mX24/M3 N_VDD_X24/M3_d N_28_X24/M3_g N_27_X24/M3_s N_VDD_X24/M2_b P_18 L=1.8e-07
+ W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06 PS=9.3e-07
mX25/M0 N_X25/6_X25/M0_d N_51_X25/M0_g N_VSS_X25/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07 PS=7.88e-06
mX25/M1 N_31_X25/M1_d N_29_X25/M1_g N_X25/6_X25/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06 PS=9.3e-07
mX25/M2 N_31_X25/M2_d N_51_X25/M2_g N_VDD_X25/M2_s N_VDD_X25/M2_b P_18 L=1.8e-07
+ W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07 PS=7.88e-06
mX25/M3 N_VDD_X25/M3_d N_29_X25/M3_g N_31_X25/M3_s N_VDD_X25/M2_b P_18 L=1.8e-07
+ W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06 PS=9.3e-07
mX26/M0 N_X26/6_X26/M0_d N_28_X26/M0_g N_VSS_X26/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07 PS=7.88e-06
mX26/M1 N_30_X26/M1_d N_STATE0_X26/M1_g N_X26/6_X26/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06 PS=9.3e-07
mX26/M2 N_30_X26/M2_d N_28_X26/M2_g N_VDD_X26/M2_s N_VDD_X26/M2_b P_18 L=1.8e-07
+ W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07 PS=7.88e-06
mX26/M3 N_VDD_X26/M3_d N_STATE0_X26/M3_g N_30_X26/M3_s N_VDD_X26/M2_b P_18
+ L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06 PS=9.3e-07
mX27/M0 N_X27/6_X27/M0_d N_STATE0_X27/M0_g N_VSS_X27/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07 PS=7.88e-06
mX27/M1 N_32_X27/M1_d N_STATE1_X27/M1_g N_X27/6_X27/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06 PS=9.3e-07
mX27/M2 N_32_X27/M2_d N_STATE0_X27/M2_g N_VDD_X27/M2_s N_VDD_X27/M2_b P_18
+ L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07 PS=7.88e-06
mX27/M3 N_VDD_X27/M3_d N_STATE1_X27/M3_g N_32_X27/M3_s N_VDD_X27/M2_b P_18
+ L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06 PS=9.3e-07
mX28/M0 N_X28/6_X28/M0_d N_STATE1_X28/M0_g N_VSS_X28/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07 PS=7.88e-06
mX28/M1 N_33_X28/M1_d N_34_X28/M1_g N_X28/6_X28/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06 PS=9.3e-07
mX28/M2 N_33_X28/M2_d N_STATE1_X28/M2_g N_VDD_X28/M2_s N_VDD_X28/M2_b P_18
+ L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07 PS=7.88e-06
mX28/M3 N_VDD_X28/M3_d N_34_X28/M3_g N_33_X28/M3_s N_VDD_X28/M2_b P_18 L=1.8e-07
+ W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06 PS=9.3e-07
mX29/M0 N_X29/6_X29/M0_d N_S1_X29/M0_g N_VSS_X29/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07 PS=7.88e-06
mX29/M1 N_52_X29/M1_d N_STORE_X29/M1_g N_X29/6_X29/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06 PS=9.3e-07
mX29/M2 N_52_X29/M2_d N_S1_X29/M2_g N_VDD_X29/M2_s N_VDD_X29/M2_b P_18 L=1.8e-07
+ W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07 PS=7.88e-06
mX29/M3 N_VDD_X29/M3_d N_STORE_X29/M3_g N_52_X29/M3_s N_VDD_X29/M2_b P_18
+ L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06 PS=9.3e-07
mX30/X0/M0 N_X30/X0/6_X30/X0/M0_d N_7_X30/X0/M0_g N_VSS_X30/X0/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X0/M1 N_X30/10_X30/X0/M1_d N_INIT0_X30/X0/M1_g N_X30/X0/6_X30/X0/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX30/X0/M2 N_X30/10_X30/X0/M2_d N_7_X30/X0/M2_g N_VDD_X30/X0/M2_s
+ N_VDD_X30/X0/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X0/M3 N_VDD_X30/X0/M3_d N_INIT0_X30/X0/M3_g N_X30/10_X30/X0/M3_s
+ N_VDD_X30/X0/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX30/X1/M0 N_X30/X1/6_X30/X1/M0_d N_X30/12_X30/X1/M0_g N_VSS_X30/X1/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X1/M1 N_37_X30/X1/M1_d N_X30/9_X30/X1/M1_g N_X30/X1/6_X30/X1/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX30/X1/M2 N_37_X30/X1/M2_d N_X30/12_X30/X1/M2_g N_VDD_X30/X1/M2_s
+ N_VDD_X30/X1/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X1/M3 N_VDD_X30/X1/M3_d N_X30/9_X30/X1/M3_g N_37_X30/X1/M3_s
+ N_VDD_X30/X1/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX30/X2/M0 N_X30/X2/6_X30/X2/M0_d N_X30/10_X30/X2/M0_g N_VSS_X30/X2/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X2/M1 N_38_X30/X2/M1_d N_X30/8_X30/X2/M1_g N_X30/X2/6_X30/X2/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX30/X2/M2 N_38_X30/X2/M2_d N_X30/10_X30/X2/M2_g N_VDD_X30/X2/M2_s
+ N_VDD_X30/X2/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X2/M3 N_VDD_X30/X2/M3_d N_X30/8_X30/X2/M3_g N_38_X30/X2/M3_s
+ N_VDD_X30/X2/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX30/X3/M0 N_X30/X3/6_X30/X3/M0_d N_X30/10_X30/X3/M0_g N_VSS_X30/X3/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X3/M1 N_X30/13_X30/X3/M1_d N_7_X30/X3/M1_g N_X30/X3/6_X30/X3/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX30/X3/M2 N_X30/13_X30/X3/M2_d N_X30/10_X30/X3/M2_g N_VDD_X30/X3/M2_s
+ N_VDD_X30/X3/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X3/M3 N_VDD_X30/X3/M3_d N_7_X30/X3/M3_g N_X30/13_X30/X3/M3_s
+ N_VDD_X30/X3/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX30/X4/M0 N_X30/X4/6_X30/X4/M0_d N_X30/10_X30/X4/M0_g N_VSS_X30/X4/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X4/M1 N_X30/11_X30/X4/M1_d N_INIT0_X30/X4/M1_g N_X30/X4/6_X30/X4/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX30/X4/M2 N_X30/11_X30/X4/M2_d N_X30/10_X30/X4/M2_g N_VDD_X30/X4/M2_s
+ N_VDD_X30/X4/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X4/M3 N_VDD_X30/X4/M3_d N_INIT0_X30/X4/M3_g N_X30/11_X30/X4/M3_s
+ N_VDD_X30/X4/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX30/X5/M0 N_X30/X5/6_X30/X5/M0_d N_X30/13_X30/X5/M0_g N_VSS_X30/X5/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X5/M1 N_X30/14_X30/X5/M1_d N_X30/11_X30/X5/M1_g N_X30/X5/6_X30/X5/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX30/X5/M2 N_X30/14_X30/X5/M2_d N_X30/13_X30/X5/M2_g N_VDD_X30/X5/M2_s
+ N_VDD_X30/X5/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X5/M3 N_VDD_X30/X5/M3_d N_X30/11_X30/X5/M3_g N_X30/14_X30/X5/M3_s
+ N_VDD_X30/X5/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX30/X6/M0 N_X30/X6/6_X30/X6/M0_d N_X30/14_X30/X6/M0_g N_VSS_X30/X6/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X6/M1 N_X30/8_X30/X6/M1_d N_VSS_X30/X6/M1_g N_X30/X6/6_X30/X6/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX30/X6/M2 N_X30/8_X30/X6/M2_d N_X30/14_X30/X6/M2_g N_VDD_X30/X6/M2_s
+ N_VDD_X30/X6/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X6/M3 N_VDD_X30/X6/M3_d N_VSS_X30/X6/M3_g N_X30/8_X30/X6/M3_s
+ N_VDD_X30/X6/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX30/X7/M0 N_X30/X7/6_X30/X7/M0_d N_X30/14_X30/X7/M0_g N_VSS_X30/X7/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X7/M1 N_X30/12_X30/X7/M1_d N_X30/8_X30/X7/M1_g N_X30/X7/6_X30/X7/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX30/X7/M2 N_X30/12_X30/X7/M2_d N_X30/14_X30/X7/M2_g N_VDD_X30/X7/M2_s
+ N_VDD_X30/X7/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X7/M3 N_VDD_X30/X7/M3_d N_X30/8_X30/X7/M3_g N_X30/12_X30/X7/M3_s
+ N_VDD_X30/X7/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX30/X8/M0 N_X30/X8/6_X30/X8/M0_d N_VSS_X30/X8/M0_g N_VSS_X30/X8/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X8/M1 N_X30/9_X30/X8/M1_d N_X30/8_X30/X8/M1_g N_X30/X8/6_X30/X8/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX30/X8/M2 N_X30/9_X30/X8/M2_d N_VSS_X30/X8/M2_g N_VDD_X30/X8/M2_s
+ N_VDD_X30/X8/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX30/X8/M3 N_VDD_X30/X8/M3_d N_X30/8_X30/X8/M3_g N_X30/9_X30/X8/M3_s
+ N_VDD_X30/X8/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X0/M0 N_X31/X0/6_X31/X0/M0_d N_23_X31/X0/M0_g N_VSS_X31/X0/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X0/M1 N_X31/10_X31/X0/M1_d N_INIT1_X31/X0/M1_g N_X31/X0/6_X31/X0/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X0/M2 N_X31/10_X31/X0/M2_d N_23_X31/X0/M2_g N_VDD_X31/X0/M2_s
+ N_VDD_X31/X0/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X0/M3 N_VDD_X31/X0/M3_d N_INIT1_X31/X0/M3_g N_X31/10_X31/X0/M3_s
+ N_VDD_X31/X0/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X1/M0 N_X31/X1/6_X31/X1/M0_d N_X31/12_X31/X1/M0_g N_VSS_X31/X1/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X1/M1 N_21_X31/X1/M1_d N_X31/9_X31/X1/M1_g N_X31/X1/6_X31/X1/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X1/M2 N_21_X31/X1/M2_d N_X31/12_X31/X1/M2_g N_VDD_X31/X1/M2_s
+ N_VDD_X31/X1/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X1/M3 N_VDD_X31/X1/M3_d N_X31/9_X31/X1/M3_g N_21_X31/X1/M3_s
+ N_VDD_X31/X1/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X2/M0 N_X31/X2/6_X31/X2/M0_d N_X31/10_X31/X2/M0_g N_VSS_X31/X2/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X2/M1 N_39_X31/X2/M1_d N_X31/8_X31/X2/M1_g N_X31/X2/6_X31/X2/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X2/M2 N_39_X31/X2/M2_d N_X31/10_X31/X2/M2_g N_VDD_X31/X2/M2_s
+ N_VDD_X31/X2/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X2/M3 N_VDD_X31/X2/M3_d N_X31/8_X31/X2/M3_g N_39_X31/X2/M3_s
+ N_VDD_X31/X2/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X3/M0 N_X31/X3/6_X31/X3/M0_d N_X31/10_X31/X3/M0_g N_VSS_X31/X3/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X3/M1 N_X31/13_X31/X3/M1_d N_23_X31/X3/M1_g N_X31/X3/6_X31/X3/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X3/M2 N_X31/13_X31/X3/M2_d N_X31/10_X31/X3/M2_g N_VDD_X31/X3/M2_s
+ N_VDD_X31/X3/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X3/M3 N_VDD_X31/X3/M3_d N_23_X31/X3/M3_g N_X31/13_X31/X3/M3_s
+ N_VDD_X31/X3/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X4/M0 N_X31/X4/6_X31/X4/M0_d N_X31/10_X31/X4/M0_g N_VSS_X31/X4/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X4/M1 N_X31/11_X31/X4/M1_d N_INIT1_X31/X4/M1_g N_X31/X4/6_X31/X4/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X4/M2 N_X31/11_X31/X4/M2_d N_X31/10_X31/X4/M2_g N_VDD_X31/X4/M2_s
+ N_VDD_X31/X4/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X4/M3 N_VDD_X31/X4/M3_d N_INIT1_X31/X4/M3_g N_X31/11_X31/X4/M3_s
+ N_VDD_X31/X4/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X5/M0 N_X31/X5/6_X31/X5/M0_d N_X31/13_X31/X5/M0_g N_VSS_X31/X5/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X5/M1 N_X31/14_X31/X5/M1_d N_X31/11_X31/X5/M1_g N_X31/X5/6_X31/X5/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X5/M2 N_X31/14_X31/X5/M2_d N_X31/13_X31/X5/M2_g N_VDD_X31/X5/M2_s
+ N_VDD_X31/X5/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X5/M3 N_VDD_X31/X5/M3_d N_X31/11_X31/X5/M3_g N_X31/14_X31/X5/M3_s
+ N_VDD_X31/X5/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X6/M0 N_X31/X6/6_X31/X6/M0_d N_X31/14_X31/X6/M0_g N_VSS_X31/X6/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X6/M1 N_X31/8_X31/X6/M1_d N_38_X31/X6/M1_g N_X31/X6/6_X31/X6/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X6/M2 N_X31/8_X31/X6/M2_d N_X31/14_X31/X6/M2_g N_VDD_X31/X6/M2_s
+ N_VDD_X31/X6/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X6/M3 N_VDD_X31/X6/M3_d N_38_X31/X6/M3_g N_X31/8_X31/X6/M3_s
+ N_VDD_X31/X6/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X7/M0 N_X31/X7/6_X31/X7/M0_d N_X31/14_X31/X7/M0_g N_VSS_X31/X7/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X7/M1 N_X31/12_X31/X7/M1_d N_X31/8_X31/X7/M1_g N_X31/X7/6_X31/X7/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X7/M2 N_X31/12_X31/X7/M2_d N_X31/14_X31/X7/M2_g N_VDD_X31/X7/M2_s
+ N_VDD_X31/X7/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X7/M3 N_VDD_X31/X7/M3_d N_X31/8_X31/X7/M3_g N_X31/12_X31/X7/M3_s
+ N_VDD_X31/X7/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X8/M0 N_X31/X8/6_X31/X8/M0_d N_38_X31/X8/M0_g N_VSS_X31/X8/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X8/M1 N_X31/9_X31/X8/M1_d N_X31/8_X31/X8/M1_g N_X31/X8/6_X31/X8/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX31/X8/M2 N_X31/9_X31/X8/M2_d N_38_X31/X8/M2_g N_VDD_X31/X8/M2_s
+ N_VDD_X31/X8/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX31/X8/M3 N_VDD_X31/X8/M3_d N_X31/8_X31/X8/M3_g N_X31/9_X31/X8/M3_s
+ N_VDD_X31/X8/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X0/M0 N_X32/X0/6_X32/X0/M0_d N_20_X32/X0/M0_g N_VSS_X32/X0/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X0/M1 N_X32/10_X32/X0/M1_d N_INIT2_X32/X0/M1_g N_X32/X0/6_X32/X0/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X0/M2 N_X32/10_X32/X0/M2_d N_20_X32/X0/M2_g N_VDD_X32/X0/M2_s
+ N_VDD_X32/X0/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X0/M3 N_VDD_X32/X0/M3_d N_INIT2_X32/X0/M3_g N_X32/10_X32/X0/M3_s
+ N_VDD_X32/X0/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X1/M0 N_X32/X1/6_X32/X1/M0_d N_X32/12_X32/X1/M0_g N_VSS_X32/X1/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X1/M1 N_22_X32/X1/M1_d N_X32/9_X32/X1/M1_g N_X32/X1/6_X32/X1/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X1/M2 N_22_X32/X1/M2_d N_X32/12_X32/X1/M2_g N_VDD_X32/X1/M2_s
+ N_VDD_X32/X1/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X1/M3 N_VDD_X32/X1/M3_d N_X32/9_X32/X1/M3_g N_22_X32/X1/M3_s
+ N_VDD_X32/X1/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X2/M0 N_X32/X2/6_X32/X2/M0_d N_X32/10_X32/X2/M0_g N_VSS_X32/X2/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X2/M1 N_40_X32/X2/M1_d N_X32/8_X32/X2/M1_g N_X32/X2/6_X32/X2/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X2/M2 N_40_X32/X2/M2_d N_X32/10_X32/X2/M2_g N_VDD_X32/X2/M2_s
+ N_VDD_X32/X2/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X2/M3 N_VDD_X32/X2/M3_d N_X32/8_X32/X2/M3_g N_40_X32/X2/M3_s
+ N_VDD_X32/X2/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X3/M0 N_X32/X3/6_X32/X3/M0_d N_X32/10_X32/X3/M0_g N_VSS_X32/X3/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X3/M1 N_X32/13_X32/X3/M1_d N_20_X32/X3/M1_g N_X32/X3/6_X32/X3/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X3/M2 N_X32/13_X32/X3/M2_d N_X32/10_X32/X3/M2_g N_VDD_X32/X3/M2_s
+ N_VDD_X32/X3/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X3/M3 N_VDD_X32/X3/M3_d N_20_X32/X3/M3_g N_X32/13_X32/X3/M3_s
+ N_VDD_X32/X3/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X4/M0 N_X32/X4/6_X32/X4/M0_d N_X32/10_X32/X4/M0_g N_VSS_X32/X4/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X4/M1 N_X32/11_X32/X4/M1_d N_INIT2_X32/X4/M1_g N_X32/X4/6_X32/X4/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X4/M2 N_X32/11_X32/X4/M2_d N_X32/10_X32/X4/M2_g N_VDD_X32/X4/M2_s
+ N_VDD_X32/X4/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X4/M3 N_VDD_X32/X4/M3_d N_INIT2_X32/X4/M3_g N_X32/11_X32/X4/M3_s
+ N_VDD_X32/X4/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X5/M0 N_X32/X5/6_X32/X5/M0_d N_X32/13_X32/X5/M0_g N_VSS_X32/X5/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X5/M1 N_X32/14_X32/X5/M1_d N_X32/11_X32/X5/M1_g N_X32/X5/6_X32/X5/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X5/M2 N_X32/14_X32/X5/M2_d N_X32/13_X32/X5/M2_g N_VDD_X32/X5/M2_s
+ N_VDD_X32/X5/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X5/M3 N_VDD_X32/X5/M3_d N_X32/11_X32/X5/M3_g N_X32/14_X32/X5/M3_s
+ N_VDD_X32/X5/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X6/M0 N_X32/X6/6_X32/X6/M0_d N_X32/14_X32/X6/M0_g N_VSS_X32/X6/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X6/M1 N_X32/8_X32/X6/M1_d N_39_X32/X6/M1_g N_X32/X6/6_X32/X6/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X6/M2 N_X32/8_X32/X6/M2_d N_X32/14_X32/X6/M2_g N_VDD_X32/X6/M2_s
+ N_VDD_X32/X6/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X6/M3 N_VDD_X32/X6/M3_d N_39_X32/X6/M3_g N_X32/8_X32/X6/M3_s
+ N_VDD_X32/X6/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X7/M0 N_X32/X7/6_X32/X7/M0_d N_X32/14_X32/X7/M0_g N_VSS_X32/X7/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X7/M1 N_X32/12_X32/X7/M1_d N_X32/8_X32/X7/M1_g N_X32/X7/6_X32/X7/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X7/M2 N_X32/12_X32/X7/M2_d N_X32/14_X32/X7/M2_g N_VDD_X32/X7/M2_s
+ N_VDD_X32/X7/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X7/M3 N_VDD_X32/X7/M3_d N_X32/8_X32/X7/M3_g N_X32/12_X32/X7/M3_s
+ N_VDD_X32/X7/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X8/M0 N_X32/X8/6_X32/X8/M0_d N_39_X32/X8/M0_g N_VSS_X32/X8/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X8/M1 N_X32/9_X32/X8/M1_d N_X32/8_X32/X8/M1_g N_X32/X8/6_X32/X8/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX32/X8/M2 N_X32/9_X32/X8/M2_d N_39_X32/X8/M2_g N_VDD_X32/X8/M2_s
+ N_VDD_X32/X8/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX32/X8/M3 N_VDD_X32/X8/M3_d N_X32/8_X32/X8/M3_g N_X32/9_X32/X8/M3_s
+ N_VDD_X32/X8/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X0/M0 N_X33/X0/6_X33/X0/M0_d N_14_X33/X0/M0_g N_VSS_X33/X0/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X0/M1 N_X33/10_X33/X0/M1_d N_INIT3_X33/X0/M1_g N_X33/X0/6_X33/X0/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X0/M2 N_X33/10_X33/X0/M2_d N_14_X33/X0/M2_g N_VDD_X33/X0/M2_s
+ N_VDD_X33/X0/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X0/M3 N_VDD_X33/X0/M3_d N_INIT3_X33/X0/M3_g N_X33/10_X33/X0/M3_s
+ N_VDD_X33/X0/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X1/M0 N_X33/X1/6_X33/X1/M0_d N_X33/12_X33/X1/M0_g N_VSS_X33/X1/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X1/M1 N_19_X33/X1/M1_d N_X33/9_X33/X1/M1_g N_X33/X1/6_X33/X1/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X1/M2 N_19_X33/X1/M2_d N_X33/12_X33/X1/M2_g N_VDD_X33/X1/M2_s
+ N_VDD_X33/X1/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X1/M3 N_VDD_X33/X1/M3_d N_X33/9_X33/X1/M3_g N_19_X33/X1/M3_s
+ N_VDD_X33/X1/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X2/M0 N_X33/X2/6_X33/X2/M0_d N_X33/10_X33/X2/M0_g N_VSS_X33/X2/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X2/M1 N_53_X33/X2/M1_d N_X33/8_X33/X2/M1_g N_X33/X2/6_X33/X2/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X2/M2 N_53_X33/X2/M2_d N_X33/10_X33/X2/M2_g N_VDD_X33/X2/M2_s
+ N_VDD_X33/X2/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X2/M3 N_VDD_X33/X2/M3_d N_X33/8_X33/X2/M3_g N_53_X33/X2/M3_s
+ N_VDD_X33/X2/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X3/M0 N_X33/X3/6_X33/X3/M0_d N_X33/10_X33/X3/M0_g N_VSS_X33/X3/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X3/M1 N_X33/13_X33/X3/M1_d N_14_X33/X3/M1_g N_X33/X3/6_X33/X3/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X3/M2 N_X33/13_X33/X3/M2_d N_X33/10_X33/X3/M2_g N_VDD_X33/X3/M2_s
+ N_VDD_X33/X3/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X3/M3 N_VDD_X33/X3/M3_d N_14_X33/X3/M3_g N_X33/13_X33/X3/M3_s
+ N_VDD_X33/X3/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X4/M0 N_X33/X4/6_X33/X4/M0_d N_X33/10_X33/X4/M0_g N_VSS_X33/X4/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X4/M1 N_X33/11_X33/X4/M1_d N_INIT3_X33/X4/M1_g N_X33/X4/6_X33/X4/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X4/M2 N_X33/11_X33/X4/M2_d N_X33/10_X33/X4/M2_g N_VDD_X33/X4/M2_s
+ N_VDD_X33/X4/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X4/M3 N_VDD_X33/X4/M3_d N_INIT3_X33/X4/M3_g N_X33/11_X33/X4/M3_s
+ N_VDD_X33/X4/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X5/M0 N_X33/X5/6_X33/X5/M0_d N_X33/13_X33/X5/M0_g N_VSS_X33/X5/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X5/M1 N_X33/14_X33/X5/M1_d N_X33/11_X33/X5/M1_g N_X33/X5/6_X33/X5/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X5/M2 N_X33/14_X33/X5/M2_d N_X33/13_X33/X5/M2_g N_VDD_X33/X5/M2_s
+ N_VDD_X33/X5/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X5/M3 N_VDD_X33/X5/M3_d N_X33/11_X33/X5/M3_g N_X33/14_X33/X5/M3_s
+ N_VDD_X33/X5/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X6/M0 N_X33/X6/6_X33/X6/M0_d N_X33/14_X33/X6/M0_g N_VSS_X33/X6/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X6/M1 N_X33/8_X33/X6/M1_d N_40_X33/X6/M1_g N_X33/X6/6_X33/X6/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X6/M2 N_X33/8_X33/X6/M2_d N_X33/14_X33/X6/M2_g N_VDD_X33/X6/M2_s
+ N_VDD_X33/X6/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X6/M3 N_VDD_X33/X6/M3_d N_40_X33/X6/M3_g N_X33/8_X33/X6/M3_s
+ N_VDD_X33/X6/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X7/M0 N_X33/X7/6_X33/X7/M0_d N_X33/14_X33/X7/M0_g N_VSS_X33/X7/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X7/M1 N_X33/12_X33/X7/M1_d N_X33/8_X33/X7/M1_g N_X33/X7/6_X33/X7/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X7/M2 N_X33/12_X33/X7/M2_d N_X33/14_X33/X7/M2_g N_VDD_X33/X7/M2_s
+ N_VDD_X33/X7/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X7/M3 N_VDD_X33/X7/M3_d N_X33/8_X33/X7/M3_g N_X33/12_X33/X7/M3_s
+ N_VDD_X33/X7/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X8/M0 N_X33/X8/6_X33/X8/M0_d N_40_X33/X8/M0_g N_VSS_X33/X8/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X8/M1 N_X33/9_X33/X8/M1_d N_X33/8_X33/X8/M1_g N_X33/X8/6_X33/X8/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX33/X8/M2 N_X33/9_X33/X8/M2_d N_40_X33/X8/M2_g N_VDD_X33/X8/M2_s
+ N_VDD_X33/X8/M2_b P_18 L=1.8e-07 W=6e-06 AD=2.79e-12 AS=5.64e-12 PD=9.3e-07
+ PS=7.88e-06
mX33/X8/M3 N_VDD_X33/X8/M3_d N_X33/8_X33/X8/M3_g N_X33/9_X33/X8/M3_s
+ N_VDD_X33/X8/M2_b P_18 L=1.8e-07 W=6e-06 AD=5.4e-12 AS=2.79e-12 PD=7.8e-06
+ PS=9.3e-07
mX34/M0 N_X34/8_X34/M0_d N_35_X34/M0_g N_VSS_X34/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.59e-12 AS=1.86e-12 PD=4.06e-06 PS=4.24e-06
mX34/M1 N_X34/10_X34/M1_d N_X34/8_X34/M1_g N_VSS_X34/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=7.95e-13 AS=1.5e-12 PD=5.3e-07 PS=4e-06
mX34/M2 N_X34/7_X34/M2_d N_VSS_X34/M2_g N_X34/10_X34/M2_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.59e-12 AS=7.95e-13 PD=4.06e-06 PS=5.3e-07
mX34/M3 N_X34/11_X34/M3_d N_35_X34/M3_g N_VSS_X34/M3_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=8.55e-13 AS=1.5e-12 PD=5.7e-07 PS=4e-06
mX34/M4 N_X34/9_X34/M4_d N_M3_X34/M4_g N_X34/11_X34/M4_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.62e-12 AS=8.55e-13 PD=4.08e-06 PS=5.7e-07
mX34/M5 N_X34/12_X34/M5_d N_X34/9_X34/M5_g N_VSS_X34/M5_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.86e-12 PD=9.8e-07 PS=4.24e-06
mX34/M6 N_16_X34/M6_d N_X34/7_X34/M6_g N_X34/12_X34/M6_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.62e-12 AS=1.47e-12 PD=4.08e-06 PS=9.8e-07
mX34/M7 N_X34/8_X34/M7_d N_35_X34/M7_g N_VDD_X34/M7_s N_VDD_X34/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=5.456e-12 PD=9.86e-06 PS=1.004e-05
mX34/M8 N_X34/7_X34/M8_d N_X34/8_X34/M8_g N_VDD_X34/M8_s N_VDD_X34/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=2.332e-12 AS=4.4e-12 PD=5.3e-07 PS=9.8e-06
mX34/M9 N_VDD_X34/M9_d N_VSS_X34/M9_g N_X34/7_X34/M9_s N_VDD_X34/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=2.332e-12 PD=9.86e-06 PS=5.3e-07
mX34/M10 N_X34/9_X34/M10_d N_35_X34/M10_g N_VDD_X34/M10_s N_VDD_X34/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=2.508e-12 AS=4.4e-12 PD=5.7e-07 PS=9.8e-06
mX34/M11 N_VDD_X34/M11_d N_M3_X34/M11_g N_X34/9_X34/M11_s N_VDD_X34/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=5.192e-12 AS=2.508e-12 PD=9.98e-06 PS=5.7e-07
mX34/M12 N_16_X34/M12_d N_X34/9_X34/M12_g N_VDD_X34/M12_s N_VDD_X34/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=4.312e-12 AS=5.016e-12 PD=9.8e-07 PS=9.94e-06
mX34/M13 N_VDD_X34/M13_d N_X34/7_X34/M13_g N_16_X34/M13_s N_VDD_X34/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=4.312e-12 PD=9.86e-06 PS=9.8e-07
mX35/M0 N_X35/8_X35/M0_d N_35_X35/M0_g N_VSS_X35/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.59e-12 AS=1.86e-12 PD=4.06e-06 PS=4.24e-06
mX35/M1 N_X35/10_X35/M1_d N_X35/8_X35/M1_g N_VSS_X35/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=7.95e-13 AS=1.5e-12 PD=5.3e-07 PS=4e-06
mX35/M2 N_X35/7_X35/M2_d N_VSS_X35/M2_g N_X35/10_X35/M2_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.59e-12 AS=7.95e-13 PD=4.06e-06 PS=5.3e-07
mX35/M3 N_X35/11_X35/M3_d N_35_X35/M3_g N_VSS_X35/M3_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=8.55e-13 AS=1.5e-12 PD=5.7e-07 PS=4e-06
mX35/M4 N_X35/9_X35/M4_d N_M1_X35/M4_g N_X35/11_X35/M4_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.62e-12 AS=8.55e-13 PD=4.08e-06 PS=5.7e-07
mX35/M5 N_X35/12_X35/M5_d N_X35/9_X35/M5_g N_VSS_X35/M5_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.86e-12 PD=9.8e-07 PS=4.24e-06
mX35/M6 N_36_X35/M6_d N_X35/7_X35/M6_g N_X35/12_X35/M6_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.62e-12 AS=1.47e-12 PD=4.08e-06 PS=9.8e-07
mX35/M7 N_X35/8_X35/M7_d N_35_X35/M7_g N_VDD_X35/M7_s N_VDD_X35/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=5.456e-12 PD=9.86e-06 PS=1.004e-05
mX35/M8 N_X35/7_X35/M8_d N_X35/8_X35/M8_g N_VDD_X35/M8_s N_VDD_X35/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=2.332e-12 AS=4.4e-12 PD=5.3e-07 PS=9.8e-06
mX35/M9 N_VDD_X35/M9_d N_VSS_X35/M9_g N_X35/7_X35/M9_s N_VDD_X35/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=2.332e-12 PD=9.86e-06 PS=5.3e-07
mX35/M10 N_X35/9_X35/M10_d N_35_X35/M10_g N_VDD_X35/M10_s N_VDD_X35/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=2.508e-12 AS=4.4e-12 PD=5.7e-07 PS=9.8e-06
mX35/M11 N_VDD_X35/M11_d N_M1_X35/M11_g N_X35/9_X35/M11_s N_VDD_X35/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=5.192e-12 AS=2.508e-12 PD=9.98e-06 PS=5.7e-07
mX35/M12 N_36_X35/M12_d N_X35/9_X35/M12_g N_VDD_X35/M12_s N_VDD_X35/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=4.312e-12 AS=5.016e-12 PD=9.8e-07 PS=9.94e-06
mX35/M13 N_VDD_X35/M13_d N_X35/7_X35/M13_g N_36_X35/M13_s N_VDD_X35/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=4.312e-12 PD=9.86e-06 PS=9.8e-07
mX36/M0 N_X36/8_X36/M0_d N_35_X36/M0_g N_VSS_X36/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.59e-12 AS=1.86e-12 PD=4.06e-06 PS=4.24e-06
mX36/M1 N_X36/10_X36/M1_d N_X36/8_X36/M1_g N_VSS_X36/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=7.95e-13 AS=1.5e-12 PD=5.3e-07 PS=4e-06
mX36/M2 N_X36/7_X36/M2_d N_VSS_X36/M2_g N_X36/10_X36/M2_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.59e-12 AS=7.95e-13 PD=4.06e-06 PS=5.3e-07
mX36/M3 N_X36/11_X36/M3_d N_35_X36/M3_g N_VSS_X36/M3_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=8.55e-13 AS=1.5e-12 PD=5.7e-07 PS=4e-06
mX36/M4 N_X36/9_X36/M4_d N_M2_X36/M4_g N_X36/11_X36/M4_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.62e-12 AS=8.55e-13 PD=4.08e-06 PS=5.7e-07
mX36/M5 N_X36/12_X36/M5_d N_X36/9_X36/M5_g N_VSS_X36/M5_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.86e-12 PD=9.8e-07 PS=4.24e-06
mX36/M6 N_18_X36/M6_d N_X36/7_X36/M6_g N_X36/12_X36/M6_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.62e-12 AS=1.47e-12 PD=4.08e-06 PS=9.8e-07
mX36/M7 N_X36/8_X36/M7_d N_35_X36/M7_g N_VDD_X36/M7_s N_VDD_X36/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=5.456e-12 PD=9.86e-06 PS=1.004e-05
mX36/M8 N_X36/7_X36/M8_d N_X36/8_X36/M8_g N_VDD_X36/M8_s N_VDD_X36/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=2.332e-12 AS=4.4e-12 PD=5.3e-07 PS=9.8e-06
mX36/M9 N_VDD_X36/M9_d N_VSS_X36/M9_g N_X36/7_X36/M9_s N_VDD_X36/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=2.332e-12 PD=9.86e-06 PS=5.3e-07
mX36/M10 N_X36/9_X36/M10_d N_35_X36/M10_g N_VDD_X36/M10_s N_VDD_X36/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=2.508e-12 AS=4.4e-12 PD=5.7e-07 PS=9.8e-06
mX36/M11 N_VDD_X36/M11_d N_M2_X36/M11_g N_X36/9_X36/M11_s N_VDD_X36/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=5.192e-12 AS=2.508e-12 PD=9.98e-06 PS=5.7e-07
mX36/M12 N_18_X36/M12_d N_X36/9_X36/M12_g N_VDD_X36/M12_s N_VDD_X36/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=4.312e-12 AS=5.016e-12 PD=9.8e-07 PS=9.94e-06
mX36/M13 N_VDD_X36/M13_d N_X36/7_X36/M13_g N_18_X36/M13_s N_VDD_X36/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=4.312e-12 PD=9.86e-06 PS=9.8e-07
mX37/M0 N_X37/8_X37/M0_d N_35_X37/M0_g N_VSS_X37/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.59e-12 AS=1.86e-12 PD=4.06e-06 PS=4.24e-06
mX37/M1 N_X37/10_X37/M1_d N_X37/8_X37/M1_g N_VSS_X37/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=7.95e-13 AS=1.5e-12 PD=5.3e-07 PS=4e-06
mX37/M2 N_X37/7_X37/M2_d N_VSS_X37/M2_g N_X37/10_X37/M2_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.59e-12 AS=7.95e-13 PD=4.06e-06 PS=5.3e-07
mX37/M3 N_X37/11_X37/M3_d N_35_X37/M3_g N_VSS_X37/M3_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=8.55e-13 AS=1.5e-12 PD=5.7e-07 PS=4e-06
mX37/M4 N_X37/9_X37/M4_d N_M0_X37/M4_g N_X37/11_X37/M4_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.62e-12 AS=8.55e-13 PD=4.08e-06 PS=5.7e-07
mX37/M5 N_X37/12_X37/M5_d N_X37/9_X37/M5_g N_VSS_X37/M5_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.86e-12 PD=9.8e-07 PS=4.24e-06
mX37/M6 N_17_X37/M6_d N_X37/7_X37/M6_g N_X37/12_X37/M6_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=1.62e-12 AS=1.47e-12 PD=4.08e-06 PS=9.8e-07
mX37/M7 N_X37/8_X37/M7_d N_35_X37/M7_g N_VDD_X37/M7_s N_VDD_X37/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=5.456e-12 PD=9.86e-06 PS=1.004e-05
mX37/M8 N_X37/7_X37/M8_d N_X37/8_X37/M8_g N_VDD_X37/M8_s N_VDD_X37/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=2.332e-12 AS=4.4e-12 PD=5.3e-07 PS=9.8e-06
mX37/M9 N_VDD_X37/M9_d N_VSS_X37/M9_g N_X37/7_X37/M9_s N_VDD_X37/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=2.332e-12 PD=9.86e-06 PS=5.3e-07
mX37/M10 N_X37/9_X37/M10_d N_35_X37/M10_g N_VDD_X37/M10_s N_VDD_X37/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=2.508e-12 AS=4.4e-12 PD=5.7e-07 PS=9.8e-06
mX37/M11 N_VDD_X37/M11_d N_M0_X37/M11_g N_X37/9_X37/M11_s N_VDD_X37/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=5.192e-12 AS=2.508e-12 PD=9.98e-06 PS=5.7e-07
mX37/M12 N_17_X37/M12_d N_X37/9_X37/M12_g N_VDD_X37/M12_s N_VDD_X37/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=4.312e-12 AS=5.016e-12 PD=9.8e-07 PS=9.94e-06
mX37/M13 N_VDD_X37/M13_d N_X37/7_X37/M13_g N_17_X37/M13_s N_VDD_X37/M7_b P_18
+ L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=4.312e-12 PD=9.86e-06 PS=9.8e-07
mX38/M0 N_X38/7_X38/M0_d N_5_X38/M0_g N_VSS_X38/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.32e-12 AS=2.72e-12 PD=5.16e-06 PS=5.36e-06
mX38/M1 N_X38/10_X38/M1_d N_CLK_X38/M1_g N_VSS_X38/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=1.28e-12 AS=3.16e-12 PD=6.4e-07 PS=5.58e-06
mX38/M2 N_X38/8_X38/M2_d N_X38/7_X38/M2_g N_X38/10_X38/M2_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.52e-12 AS=1.28e-12 PD=5.26e-06 PS=6.4e-07
mX38/M3 N_X38/11_X38/M3_d N_X38/8_X38/M3_g N_VSS_X38/M3_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=9.8e-13 AS=2.2e-12 PD=4.9e-07 PS=5.1e-06
mX38/M4 N_6_X38/M4_d N_CLK_X38/M4_g N_X38/11_X38/M4_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.08e-12 AS=9.8e-13 PD=5.04e-06 PS=4.9e-07
mX38/M5 N_STATE0_X38/M5_d N_6_X38/M5_g N_VSS_X38/M5_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.56e-12 AS=2.08e-12 PD=5.28e-06 PS=5.04e-06
mX38/M6 N_X38/9_X38/M6_d N_5_X38/M6_g N_VDD_X38/M6_s N_VDD_X38/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=2.8635e-12 AS=5.644e-12 PD=6.9e-07 PS=9.66e-06
mX38/M7 N_X38/7_X38/M7_d N_CLK_X38/M7_g N_X38/9_X38/M7_s N_VDD_X38/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.81e-12 AS=2.8635e-12 PD=9.7e-06 PS=6.9e-07
mX38/M8 N_X38/8_X38/M8_d N_CLK_X38/M8_g N_VDD_X38/M8_s N_VDD_X38/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.644e-12 AS=5.395e-12 PD=9.66e-06 PS=9.6e-06
mX38/M9 N_6_X38/M9_d N_X38/8_X38/M9_g N_VDD_X38/M9_s N_VDD_X38/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.478e-12 AS=5.063e-12 PD=9.62e-06 PS=9.52e-06
mX38/M10 N_STATE0_X38/M10_d N_6_X38/M10_g N_VDD_X38/M10_s N_VDD_X38/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.229e-12 AS=6.557e-12 PD=9.56e-06 PS=9.88e-06
mX39/M0 N_X39/7_X39/M0_d N_31_X39/M0_g N_VSS_X39/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.32e-12 AS=2.72e-12 PD=5.16e-06 PS=5.36e-06
mX39/M1 N_X39/10_X39/M1_d N_CLK_X39/M1_g N_VSS_X39/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=1.28e-12 AS=3.16e-12 PD=6.4e-07 PS=5.58e-06
mX39/M2 N_X39/8_X39/M2_d N_X39/7_X39/M2_g N_X39/10_X39/M2_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.52e-12 AS=1.28e-12 PD=5.26e-06 PS=6.4e-07
mX39/M3 N_X39/11_X39/M3_d N_X39/8_X39/M3_g N_VSS_X39/M3_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=9.8e-13 AS=2.2e-12 PD=4.9e-07 PS=5.1e-06
mX39/M4 N_11_X39/M4_d N_CLK_X39/M4_g N_X39/11_X39/M4_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.08e-12 AS=9.8e-13 PD=5.04e-06 PS=4.9e-07
mX39/M5 N_STATE1_X39/M5_d N_11_X39/M5_g N_VSS_X39/M5_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.56e-12 AS=2.08e-12 PD=5.28e-06 PS=5.04e-06
mX39/M6 N_X39/9_X39/M6_d N_31_X39/M6_g N_VDD_X39/M6_s N_VDD_X39/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=2.8635e-12 AS=5.644e-12 PD=6.9e-07 PS=9.66e-06
mX39/M7 N_X39/7_X39/M7_d N_CLK_X39/M7_g N_X39/9_X39/M7_s N_VDD_X39/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.81e-12 AS=2.8635e-12 PD=9.7e-06 PS=6.9e-07
mX39/M8 N_X39/8_X39/M8_d N_CLK_X39/M8_g N_VDD_X39/M8_s N_VDD_X39/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.644e-12 AS=5.395e-12 PD=9.66e-06 PS=9.6e-06
mX39/M9 N_11_X39/M9_d N_X39/8_X39/M9_g N_VDD_X39/M9_s N_VDD_X39/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.478e-12 AS=5.063e-12 PD=9.62e-06 PS=9.52e-06
mX39/M10 N_STATE1_X39/M10_d N_11_X39/M10_g N_VDD_X39/M10_s N_VDD_X39/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.229e-12 AS=6.557e-12 PD=9.56e-06 PS=9.88e-06
mX40/M0 N_X40/7_X40/M0_d N_21_X40/M0_g N_VSS_X40/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.32e-12 AS=2.72e-12 PD=5.16e-06 PS=5.36e-06
mX40/M1 N_X40/10_X40/M1_d N_CLK_X40/M1_g N_VSS_X40/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=1.28e-12 AS=3.16e-12 PD=6.4e-07 PS=5.58e-06
mX40/M2 N_X40/8_X40/M2_d N_X40/7_X40/M2_g N_X40/10_X40/M2_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.52e-12 AS=1.28e-12 PD=5.26e-06 PS=6.4e-07
mX40/M3 N_X40/11_X40/M3_d N_X40/8_X40/M3_g N_VSS_X40/M3_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=9.8e-13 AS=2.2e-12 PD=4.9e-07 PS=5.1e-06
mX40/M4 N_41_X40/M4_d N_CLK_X40/M4_g N_X40/11_X40/M4_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.08e-12 AS=9.8e-13 PD=5.04e-06 PS=4.9e-07
mX40/M5 N_INIT1_X40/M5_d N_41_X40/M5_g N_VSS_X40/M5_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.56e-12 AS=2.08e-12 PD=5.28e-06 PS=5.04e-06
mX40/M6 N_X40/9_X40/M6_d N_21_X40/M6_g N_VDD_X40/M6_s N_VDD_X40/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=2.8635e-12 AS=5.644e-12 PD=6.9e-07 PS=9.66e-06
mX40/M7 N_X40/7_X40/M7_d N_CLK_X40/M7_g N_X40/9_X40/M7_s N_VDD_X40/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.81e-12 AS=2.8635e-12 PD=9.7e-06 PS=6.9e-07
mX40/M8 N_X40/8_X40/M8_d N_CLK_X40/M8_g N_VDD_X40/M8_s N_VDD_X40/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.644e-12 AS=5.395e-12 PD=9.66e-06 PS=9.6e-06
mX40/M9 N_41_X40/M9_d N_X40/8_X40/M9_g N_VDD_X40/M9_s N_VDD_X40/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.478e-12 AS=5.063e-12 PD=9.62e-06 PS=9.52e-06
mX40/M10 N_INIT1_X40/M10_d N_41_X40/M10_g N_VDD_X40/M10_s N_VDD_X40/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.229e-12 AS=6.557e-12 PD=9.56e-06 PS=9.88e-06
mX41/M0 N_X41/7_X41/M0_d N_19_X41/M0_g N_VSS_X41/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.32e-12 AS=2.72e-12 PD=5.16e-06 PS=5.36e-06
mX41/M1 N_X41/10_X41/M1_d N_CLK_X41/M1_g N_VSS_X41/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=1.28e-12 AS=3.16e-12 PD=6.4e-07 PS=5.58e-06
mX41/M2 N_X41/8_X41/M2_d N_X41/7_X41/M2_g N_X41/10_X41/M2_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.52e-12 AS=1.28e-12 PD=5.26e-06 PS=6.4e-07
mX41/M3 N_X41/11_X41/M3_d N_X41/8_X41/M3_g N_VSS_X41/M3_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=9.8e-13 AS=2.2e-12 PD=4.9e-07 PS=5.1e-06
mX41/M4 N_42_X41/M4_d N_CLK_X41/M4_g N_X41/11_X41/M4_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.08e-12 AS=9.8e-13 PD=5.04e-06 PS=4.9e-07
mX41/M5 N_INIT3_X41/M5_d N_42_X41/M5_g N_VSS_X41/M5_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.56e-12 AS=2.08e-12 PD=5.28e-06 PS=5.04e-06
mX41/M6 N_X41/9_X41/M6_d N_19_X41/M6_g N_VDD_X41/M6_s N_VDD_X41/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=2.8635e-12 AS=5.644e-12 PD=6.9e-07 PS=9.66e-06
mX41/M7 N_X41/7_X41/M7_d N_CLK_X41/M7_g N_X41/9_X41/M7_s N_VDD_X41/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.81e-12 AS=2.8635e-12 PD=9.7e-06 PS=6.9e-07
mX41/M8 N_X41/8_X41/M8_d N_CLK_X41/M8_g N_VDD_X41/M8_s N_VDD_X41/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.644e-12 AS=5.395e-12 PD=9.66e-06 PS=9.6e-06
mX41/M9 N_42_X41/M9_d N_X41/8_X41/M9_g N_VDD_X41/M9_s N_VDD_X41/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.478e-12 AS=5.063e-12 PD=9.62e-06 PS=9.52e-06
mX41/M10 N_INIT3_X41/M10_d N_42_X41/M10_g N_VDD_X41/M10_s N_VDD_X41/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.229e-12 AS=6.557e-12 PD=9.56e-06 PS=9.88e-06
mX42/M0 N_X42/7_X42/M0_d N_16_X42/M0_g N_VSS_X42/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.32e-12 AS=2.72e-12 PD=5.16e-06 PS=5.36e-06
mX42/M1 N_X42/10_X42/M1_d N_CLK_X42/M1_g N_VSS_X42/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=1.28e-12 AS=3.16e-12 PD=6.4e-07 PS=5.58e-06
mX42/M2 N_X42/8_X42/M2_d N_X42/7_X42/M2_g N_X42/10_X42/M2_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.52e-12 AS=1.28e-12 PD=5.26e-06 PS=6.4e-07
mX42/M3 N_X42/11_X42/M3_d N_X42/8_X42/M3_g N_VSS_X42/M3_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=9.8e-13 AS=2.2e-12 PD=4.9e-07 PS=5.1e-06
mX42/M4 N_43_X42/M4_d N_CLK_X42/M4_g N_X42/11_X42/M4_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.08e-12 AS=9.8e-13 PD=5.04e-06 PS=4.9e-07
mX42/M5 N_14_X42/M5_d N_43_X42/M5_g N_VSS_X42/M5_s N_VSS_X24/M0_b N_18 L=1.8e-07
+ W=4e-06 AD=2.56e-12 AS=2.08e-12 PD=5.28e-06 PS=5.04e-06
mX42/M6 N_X42/9_X42/M6_d N_16_X42/M6_g N_VDD_X42/M6_s N_VDD_X42/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=2.8635e-12 AS=5.644e-12 PD=6.9e-07 PS=9.66e-06
mX42/M7 N_X42/7_X42/M7_d N_CLK_X42/M7_g N_X42/9_X42/M7_s N_VDD_X42/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.81e-12 AS=2.8635e-12 PD=9.7e-06 PS=6.9e-07
mX42/M8 N_X42/8_X42/M8_d N_CLK_X42/M8_g N_VDD_X42/M8_s N_VDD_X42/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.644e-12 AS=5.395e-12 PD=9.66e-06 PS=9.6e-06
mX42/M9 N_43_X42/M9_d N_X42/8_X42/M9_g N_VDD_X42/M9_s N_VDD_X42/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.478e-12 AS=5.063e-12 PD=9.62e-06 PS=9.52e-06
mX42/M10 N_14_X42/M10_d N_43_X42/M10_g N_VDD_X42/M10_s N_VDD_X42/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.229e-12 AS=6.557e-12 PD=9.56e-06 PS=9.88e-06
mX43/M0 N_X43/7_X43/M0_d N_36_X43/M0_g N_VSS_X43/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.32e-12 AS=2.72e-12 PD=5.16e-06 PS=5.36e-06
mX43/M1 N_X43/10_X43/M1_d N_CLK_X43/M1_g N_VSS_X43/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=1.28e-12 AS=3.16e-12 PD=6.4e-07 PS=5.58e-06
mX43/M2 N_X43/8_X43/M2_d N_X43/7_X43/M2_g N_X43/10_X43/M2_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.52e-12 AS=1.28e-12 PD=5.26e-06 PS=6.4e-07
mX43/M3 N_X43/11_X43/M3_d N_X43/8_X43/M3_g N_VSS_X43/M3_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=9.8e-13 AS=2.2e-12 PD=4.9e-07 PS=5.1e-06
mX43/M4 N_44_X43/M4_d N_CLK_X43/M4_g N_X43/11_X43/M4_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.08e-12 AS=9.8e-13 PD=5.04e-06 PS=4.9e-07
mX43/M5 N_23_X43/M5_d N_44_X43/M5_g N_VSS_X43/M5_s N_VSS_X24/M0_b N_18 L=1.8e-07
+ W=4e-06 AD=2.56e-12 AS=2.08e-12 PD=5.28e-06 PS=5.04e-06
mX43/M6 N_X43/9_X43/M6_d N_36_X43/M6_g N_VDD_X43/M6_s N_VDD_X43/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=2.8635e-12 AS=5.644e-12 PD=6.9e-07 PS=9.66e-06
mX43/M7 N_X43/7_X43/M7_d N_CLK_X43/M7_g N_X43/9_X43/M7_s N_VDD_X43/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.81e-12 AS=2.8635e-12 PD=9.7e-06 PS=6.9e-07
mX43/M8 N_X43/8_X43/M8_d N_CLK_X43/M8_g N_VDD_X43/M8_s N_VDD_X43/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.644e-12 AS=5.395e-12 PD=9.66e-06 PS=9.6e-06
mX43/M9 N_44_X43/M9_d N_X43/8_X43/M9_g N_VDD_X43/M9_s N_VDD_X43/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.478e-12 AS=5.063e-12 PD=9.62e-06 PS=9.52e-06
mX43/M10 N_23_X43/M10_d N_44_X43/M10_g N_VDD_X43/M10_s N_VDD_X43/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.229e-12 AS=6.557e-12 PD=9.56e-06 PS=9.88e-06
mX44/M0 N_X44/7_X44/M0_d N_22_X44/M0_g N_VSS_X44/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.32e-12 AS=2.72e-12 PD=5.16e-06 PS=5.36e-06
mX44/M1 N_X44/10_X44/M1_d N_CLK_X44/M1_g N_VSS_X44/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=1.28e-12 AS=3.16e-12 PD=6.4e-07 PS=5.58e-06
mX44/M2 N_X44/8_X44/M2_d N_X44/7_X44/M2_g N_X44/10_X44/M2_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.52e-12 AS=1.28e-12 PD=5.26e-06 PS=6.4e-07
mX44/M3 N_X44/11_X44/M3_d N_X44/8_X44/M3_g N_VSS_X44/M3_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=9.8e-13 AS=2.2e-12 PD=4.9e-07 PS=5.1e-06
mX44/M4 N_45_X44/M4_d N_CLK_X44/M4_g N_X44/11_X44/M4_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.08e-12 AS=9.8e-13 PD=5.04e-06 PS=4.9e-07
mX44/M5 N_INIT2_X44/M5_d N_45_X44/M5_g N_VSS_X44/M5_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.56e-12 AS=2.08e-12 PD=5.28e-06 PS=5.04e-06
mX44/M6 N_X44/9_X44/M6_d N_22_X44/M6_g N_VDD_X44/M6_s N_VDD_X44/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=2.8635e-12 AS=5.644e-12 PD=6.9e-07 PS=9.66e-06
mX44/M7 N_X44/7_X44/M7_d N_CLK_X44/M7_g N_X44/9_X44/M7_s N_VDD_X44/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.81e-12 AS=2.8635e-12 PD=9.7e-06 PS=6.9e-07
mX44/M8 N_X44/8_X44/M8_d N_CLK_X44/M8_g N_VDD_X44/M8_s N_VDD_X44/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.644e-12 AS=5.395e-12 PD=9.66e-06 PS=9.6e-06
mX44/M9 N_45_X44/M9_d N_X44/8_X44/M9_g N_VDD_X44/M9_s N_VDD_X44/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.478e-12 AS=5.063e-12 PD=9.62e-06 PS=9.52e-06
mX44/M10 N_INIT2_X44/M10_d N_45_X44/M10_g N_VDD_X44/M10_s N_VDD_X44/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.229e-12 AS=6.557e-12 PD=9.56e-06 PS=9.88e-06
mX45/M0 N_X45/7_X45/M0_d N_37_X45/M0_g N_VSS_X45/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.32e-12 AS=2.72e-12 PD=5.16e-06 PS=5.36e-06
mX45/M1 N_X45/10_X45/M1_d N_CLK_X45/M1_g N_VSS_X45/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=1.28e-12 AS=3.16e-12 PD=6.4e-07 PS=5.58e-06
mX45/M2 N_X45/8_X45/M2_d N_X45/7_X45/M2_g N_X45/10_X45/M2_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.52e-12 AS=1.28e-12 PD=5.26e-06 PS=6.4e-07
mX45/M3 N_X45/11_X45/M3_d N_X45/8_X45/M3_g N_VSS_X45/M3_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=9.8e-13 AS=2.2e-12 PD=4.9e-07 PS=5.1e-06
mX45/M4 N_46_X45/M4_d N_CLK_X45/M4_g N_X45/11_X45/M4_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.08e-12 AS=9.8e-13 PD=5.04e-06 PS=4.9e-07
mX45/M5 N_INIT0_X45/M5_d N_46_X45/M5_g N_VSS_X45/M5_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.56e-12 AS=2.08e-12 PD=5.28e-06 PS=5.04e-06
mX45/M6 N_X45/9_X45/M6_d N_37_X45/M6_g N_VDD_X45/M6_s N_VDD_X45/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=2.8635e-12 AS=5.644e-12 PD=6.9e-07 PS=9.66e-06
mX45/M7 N_X45/7_X45/M7_d N_CLK_X45/M7_g N_X45/9_X45/M7_s N_VDD_X45/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.81e-12 AS=2.8635e-12 PD=9.7e-06 PS=6.9e-07
mX45/M8 N_X45/8_X45/M8_d N_CLK_X45/M8_g N_VDD_X45/M8_s N_VDD_X45/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.644e-12 AS=5.395e-12 PD=9.66e-06 PS=9.6e-06
mX45/M9 N_46_X45/M9_d N_X45/8_X45/M9_g N_VDD_X45/M9_s N_VDD_X45/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.478e-12 AS=5.063e-12 PD=9.62e-06 PS=9.52e-06
mX45/M10 N_INIT0_X45/M10_d N_46_X45/M10_g N_VDD_X45/M10_s N_VDD_X45/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.229e-12 AS=6.557e-12 PD=9.56e-06 PS=9.88e-06
mX46/M0 N_X46/7_X46/M0_d N_17_X46/M0_g N_VSS_X46/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.32e-12 AS=2.72e-12 PD=5.16e-06 PS=5.36e-06
mX46/M1 N_X46/10_X46/M1_d N_CLK_X46/M1_g N_VSS_X46/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=1.28e-12 AS=3.16e-12 PD=6.4e-07 PS=5.58e-06
mX46/M2 N_X46/8_X46/M2_d N_X46/7_X46/M2_g N_X46/10_X46/M2_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.52e-12 AS=1.28e-12 PD=5.26e-06 PS=6.4e-07
mX46/M3 N_X46/11_X46/M3_d N_X46/8_X46/M3_g N_VSS_X46/M3_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=9.8e-13 AS=2.2e-12 PD=4.9e-07 PS=5.1e-06
mX46/M4 N_47_X46/M4_d N_CLK_X46/M4_g N_X46/11_X46/M4_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.08e-12 AS=9.8e-13 PD=5.04e-06 PS=4.9e-07
mX46/M5 N_7_X46/M5_d N_47_X46/M5_g N_VSS_X46/M5_s N_VSS_X24/M0_b N_18 L=1.8e-07
+ W=4e-06 AD=2.56e-12 AS=2.08e-12 PD=5.28e-06 PS=5.04e-06
mX46/M6 N_X46/9_X46/M6_d N_17_X46/M6_g N_VDD_X46/M6_s N_VDD_X46/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=2.8635e-12 AS=5.644e-12 PD=6.9e-07 PS=9.66e-06
mX46/M7 N_X46/7_X46/M7_d N_CLK_X46/M7_g N_X46/9_X46/M7_s N_VDD_X46/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.81e-12 AS=2.8635e-12 PD=9.7e-06 PS=6.9e-07
mX46/M8 N_X46/8_X46/M8_d N_CLK_X46/M8_g N_VDD_X46/M8_s N_VDD_X46/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.644e-12 AS=5.395e-12 PD=9.66e-06 PS=9.6e-06
mX46/M9 N_47_X46/M9_d N_X46/8_X46/M9_g N_VDD_X46/M9_s N_VDD_X46/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.478e-12 AS=5.063e-12 PD=9.62e-06 PS=9.52e-06
mX46/M10 N_7_X46/M10_d N_47_X46/M10_g N_VDD_X46/M10_s N_VDD_X46/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.229e-12 AS=6.557e-12 PD=9.56e-06 PS=9.88e-06
mX47/M0 N_X47/7_X47/M0_d N_18_X47/M0_g N_VSS_X47/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.32e-12 AS=2.72e-12 PD=5.16e-06 PS=5.36e-06
mX47/M1 N_X47/10_X47/M1_d N_CLK_X47/M1_g N_VSS_X47/M1_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=1.28e-12 AS=3.16e-12 PD=6.4e-07 PS=5.58e-06
mX47/M2 N_X47/8_X47/M2_d N_X47/7_X47/M2_g N_X47/10_X47/M2_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.52e-12 AS=1.28e-12 PD=5.26e-06 PS=6.4e-07
mX47/M3 N_X47/11_X47/M3_d N_X47/8_X47/M3_g N_VSS_X47/M3_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=9.8e-13 AS=2.2e-12 PD=4.9e-07 PS=5.1e-06
mX47/M4 N_48_X47/M4_d N_CLK_X47/M4_g N_X47/11_X47/M4_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=4e-06 AD=2.08e-12 AS=9.8e-13 PD=5.04e-06 PS=4.9e-07
mX47/M5 N_20_X47/M5_d N_48_X47/M5_g N_VSS_X47/M5_s N_VSS_X24/M0_b N_18 L=1.8e-07
+ W=4e-06 AD=2.56e-12 AS=2.08e-12 PD=5.28e-06 PS=5.04e-06
mX47/M6 N_X47/9_X47/M6_d N_18_X47/M6_g N_VDD_X47/M6_s N_VDD_X47/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=2.8635e-12 AS=5.644e-12 PD=6.9e-07 PS=9.66e-06
mX47/M7 N_X47/7_X47/M7_d N_CLK_X47/M7_g N_X47/9_X47/M7_s N_VDD_X47/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.81e-12 AS=2.8635e-12 PD=9.7e-06 PS=6.9e-07
mX47/M8 N_X47/8_X47/M8_d N_CLK_X47/M8_g N_VDD_X47/M8_s N_VDD_X47/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.644e-12 AS=5.395e-12 PD=9.66e-06 PS=9.6e-06
mX47/M9 N_48_X47/M9_d N_X47/8_X47/M9_g N_VDD_X47/M9_s N_VDD_X47/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.478e-12 AS=5.063e-12 PD=9.62e-06 PS=9.52e-06
mX47/M10 N_20_X47/M10_d N_48_X47/M10_g N_VDD_X47/M10_s N_VDD_X47/M6_b P_18
+ L=1.8e-07 W=8.3e-06 AD=5.229e-12 AS=6.557e-12 PD=9.56e-06 PS=9.88e-06
mX48/M0 N_50_X48/M0_d N_STORE_X48/M0_g N_VSS_X48/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=2.13e-12 AS=2.01e-12 PD=4.42e-06 PS=4.34e-06
mX48/M1 N_50_X48/M1_d N_STORE_X48/M1_g N_VDD_X48/M1_s N_VDD_X48/M1_b P_18
+ L=1.8e-07 W=6e-06 AD=4.26e-12 AS=4.02e-12 PD=7.42e-06 PS=7.34e-06
mX49/M0 N_26_X49/M0_d N_POWER_X49/M0_g N_VSS_X49/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=2.13e-12 AS=2.01e-12 PD=4.42e-06 PS=4.34e-06
mX49/M1 N_26_X49/M1_d N_POWER_X49/M1_g N_VDD_X49/M1_s N_VDD_X49/M1_b P_18
+ L=1.8e-07 W=6e-06 AD=4.26e-12 AS=4.02e-12 PD=7.42e-06 PS=7.34e-06
mX50/M0 N_S0_X50/M0_d N_27_X50/M0_g N_VSS_X50/M0_s N_VSS_X24/M0_b N_18 L=1.8e-07
+ W=3e-06 AD=2.13e-12 AS=2.01e-12 PD=4.42e-06 PS=4.34e-06
mX50/M1 N_S0_X50/M1_d N_27_X50/M1_g N_VDD_X50/M1_s N_VDD_X50/M1_b P_18 L=1.8e-07
+ W=6e-06 AD=4.26e-12 AS=4.02e-12 PD=7.42e-06 PS=7.34e-06
mX51/M0 N_28_X51/M0_d N_STATE1_X51/M0_g N_VSS_X51/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=2.13e-12 AS=2.01e-12 PD=4.42e-06 PS=4.34e-06
mX51/M1 N_28_X51/M1_d N_STATE1_X51/M1_g N_VDD_X51/M1_s N_VDD_X51/M1_b P_18
+ L=1.8e-07 W=6e-06 AD=4.26e-12 AS=4.02e-12 PD=7.42e-06 PS=7.34e-06
mX52/M0 N_S1_X52/M0_d N_30_X52/M0_g N_VSS_X52/M0_s N_VSS_X24/M0_b N_18 L=1.8e-07
+ W=3e-06 AD=2.13e-12 AS=2.01e-12 PD=4.42e-06 PS=4.34e-06
mX52/M1 N_S1_X52/M1_d N_30_X52/M1_g N_VDD_X52/M1_s N_VDD_X50/M1_b P_18 L=1.8e-07
+ W=6e-06 AD=4.26e-12 AS=4.02e-12 PD=7.42e-06 PS=7.34e-06
mX53/M0 N_S3_X53/M0_d N_32_X53/M0_g N_VSS_X53/M0_s N_VSS_X24/M0_b N_18 L=1.8e-07
+ W=3e-06 AD=2.13e-12 AS=2.01e-12 PD=4.42e-06 PS=4.34e-06
mX53/M1 N_S3_X53/M1_d N_32_X53/M1_g N_VDD_X53/M1_s N_VDD_X53/M1_b P_18 L=1.8e-07
+ W=6e-06 AD=4.26e-12 AS=4.02e-12 PD=7.42e-06 PS=7.34e-06
mX54/M0 N_34_X54/M0_d N_STATE0_X54/M0_g N_VSS_X54/M0_s N_VSS_X24/M0_b N_18
+ L=1.8e-07 W=3e-06 AD=2.13e-12 AS=2.01e-12 PD=4.42e-06 PS=4.34e-06
mX54/M1 N_34_X54/M1_d N_STATE0_X54/M1_g N_VDD_X54/M1_s N_VDD_X54/M1_b P_18
+ L=1.8e-07 W=6e-06 AD=4.26e-12 AS=4.02e-12 PD=7.42e-06 PS=7.34e-06
mX55/M0 N_S2_X55/M0_d N_33_X55/M0_g N_VSS_X55/M0_s N_VSS_X24/M0_b N_18 L=1.8e-07
+ W=3e-06 AD=2.13e-12 AS=2.01e-12 PD=4.42e-06 PS=4.34e-06
mX55/M1 N_S2_X55/M1_d N_33_X55/M1_g N_VDD_X55/M1_s N_VDD_X53/M1_b P_18 L=1.8e-07
+ W=6e-06 AD=4.26e-12 AS=4.02e-12 PD=7.42e-06 PS=7.34e-06
mX56/M0 N_35_X56/M0_d N_52_X56/M0_g N_VSS_X56/M0_s N_VSS_X24/M0_b N_18 L=1.8e-07
+ W=3e-06 AD=2.13e-12 AS=2.01e-12 PD=4.42e-06 PS=4.34e-06
mX56/M1 N_35_X56/M1_d N_52_X56/M1_g N_VDD_X56/M1_s N_VDD_X56/M1_b P_18 L=1.8e-07
+ W=6e-06 AD=4.26e-12 AS=4.02e-12 PD=7.42e-06 PS=7.34e-06
mX57/X0/M0 N_X57/X0/8_X57/X0/M0_d N_STATE0_X57/X0/M0_g N_VSS_X57/X0/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=1.86e-12 PD=4.06e-06
+ PS=4.24e-06
mX57/X0/M1 N_X57/X0/10_X57/X0/M1_d N_X57/X0/8_X57/X0/M1_g N_VSS_X57/X0/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=7.95e-13 AS=1.5e-12 PD=5.3e-07
+ PS=4e-06
mX57/X0/M2 N_X57/X0/7_X57/X0/M2_d N_VSS_X57/X0/M2_g N_X57/X0/10_X57/X0/M2_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=7.95e-13 PD=4.06e-06
+ PS=5.3e-07
mX57/X0/M3 N_X57/X0/11_X57/X0/M3_d N_STATE0_X57/X0/M3_g N_VSS_X57/X0/M3_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=8.55e-13 AS=1.5e-12 PD=5.7e-07
+ PS=4e-06
mX57/X0/M4 N_X57/X0/9_X57/X0/M4_d N_VSS_X57/X0/M4_g N_X57/X0/11_X57/X0/M4_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=8.55e-13 PD=4.08e-06
+ PS=5.7e-07
mX57/X0/M5 N_X57/X0/12_X57/X0/M5_d N_X57/X0/9_X57/X0/M5_g N_VSS_X57/X0/M5_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.86e-12 PD=9.8e-07
+ PS=4.24e-06
mX57/X0/M6 N_X57/10_X57/X0/M6_d N_X57/X0/7_X57/X0/M6_g N_X57/X0/12_X57/X0/M6_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=1.47e-12 PD=4.08e-06
+ PS=9.8e-07
mX57/X0/M7 N_X57/X0/8_X57/X0/M7_d N_STATE0_X57/X0/M7_g N_VDD_X57/X0/M7_s
+ N_VDD_X57/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=5.456e-12
+ PD=9.86e-06 PS=1.004e-05
mX57/X0/M8 N_X57/X0/7_X57/X0/M8_d N_X57/X0/8_X57/X0/M8_g N_VDD_X57/X0/M8_s
+ N_VDD_X57/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.332e-12 AS=4.4e-12 PD=5.3e-07
+ PS=9.8e-06
mX57/X0/M9 N_VDD_X57/X0/M9_d N_VSS_X57/X0/M9_g N_X57/X0/7_X57/X0/M9_s
+ N_VDD_X57/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=2.332e-12
+ PD=9.86e-06 PS=5.3e-07
mX57/X0/M10 N_X57/X0/9_X57/X0/M10_d N_STATE0_X57/X0/M10_g N_VDD_X57/X0/M10_s
+ N_VDD_X57/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.508e-12 AS=4.4e-12 PD=5.7e-07
+ PS=9.8e-06
mX57/X0/M11 N_VDD_X57/X0/M11_d N_VSS_X57/X0/M11_g N_X57/X0/9_X57/X0/M11_s
+ N_VDD_X57/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=5.192e-12 AS=2.508e-12
+ PD=9.98e-06 PS=5.7e-07
mX57/X0/M12 N_X57/10_X57/X0/M12_d N_X57/X0/9_X57/X0/M12_g N_VDD_X57/X0/M12_s
+ N_VDD_X57/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.312e-12 AS=5.016e-12
+ PD=9.8e-07 PS=9.94e-06
mX57/X0/M13 N_VDD_X57/X0/M13_d N_X57/X0/7_X57/X0/M13_g N_X57/10_X57/X0/M13_s
+ N_VDD_X57/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=4.312e-12
+ PD=9.86e-06 PS=9.8e-07
mX57/X1/M0 N_X57/X1/8_X57/X1/M0_d N_STATE1_X57/X1/M0_g N_VSS_X57/X1/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=1.86e-12 PD=4.06e-06
+ PS=4.24e-06
mX57/X1/M1 N_X57/X1/10_X57/X1/M1_d N_X57/X1/8_X57/X1/M1_g N_VSS_X57/X1/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=7.95e-13 AS=1.5e-12 PD=5.3e-07
+ PS=4e-06
mX57/X1/M2 N_X57/X1/7_X57/X1/M2_d N_X57/10_X57/X1/M2_g N_X57/X1/10_X57/X1/M2_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=7.95e-13 PD=4.06e-06
+ PS=5.3e-07
mX57/X1/M3 N_X57/X1/11_X57/X1/M3_d N_STATE1_X57/X1/M3_g N_VSS_X57/X1/M3_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=8.55e-13 AS=1.5e-12 PD=5.7e-07
+ PS=4e-06
mX57/X1/M4 N_X57/X1/9_X57/X1/M4_d N_X57/11_X57/X1/M4_g N_X57/X1/11_X57/X1/M4_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=8.55e-13 PD=4.08e-06
+ PS=5.7e-07
mX57/X1/M5 N_X57/X1/12_X57/X1/M5_d N_X57/X1/9_X57/X1/M5_g N_VSS_X57/X1/M5_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.86e-12 PD=9.8e-07
+ PS=4.24e-06
mX57/X1/M6 N_MO1_X57/X1/M6_d N_X57/X1/7_X57/X1/M6_g N_X57/X1/12_X57/X1/M6_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=1.47e-12 PD=4.08e-06
+ PS=9.8e-07
mX57/X1/M7 N_X57/X1/8_X57/X1/M7_d N_STATE1_X57/X1/M7_g N_VDD_X57/X1/M7_s
+ N_VDD_X57/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=5.456e-12
+ PD=9.86e-06 PS=1.004e-05
mX57/X1/M8 N_X57/X1/7_X57/X1/M8_d N_X57/X1/8_X57/X1/M8_g N_VDD_X57/X1/M8_s
+ N_VDD_X57/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.332e-12 AS=4.4e-12 PD=5.3e-07
+ PS=9.8e-06
mX57/X1/M9 N_VDD_X57/X1/M9_d N_X57/10_X57/X1/M9_g N_X57/X1/7_X57/X1/M9_s
+ N_VDD_X57/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=2.332e-12
+ PD=9.86e-06 PS=5.3e-07
mX57/X1/M10 N_X57/X1/9_X57/X1/M10_d N_STATE1_X57/X1/M10_g N_VDD_X57/X1/M10_s
+ N_VDD_X57/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.508e-12 AS=4.4e-12 PD=5.7e-07
+ PS=9.8e-06
mX57/X1/M11 N_VDD_X57/X1/M11_d N_X57/11_X57/X1/M11_g N_X57/X1/9_X57/X1/M11_s
+ N_VDD_X57/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=5.192e-12 AS=2.508e-12
+ PD=9.98e-06 PS=5.7e-07
mX57/X1/M12 N_MO1_X57/X1/M12_d N_X57/X1/9_X57/X1/M12_g N_VDD_X57/X1/M12_s
+ N_VDD_X57/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.312e-12 AS=5.016e-12
+ PD=9.8e-07 PS=9.94e-06
mX57/X1/M13 N_VDD_X57/X1/M13_d N_X57/X1/7_X57/X1/M13_g N_MO1_X57/X1/M13_s
+ N_VDD_X57/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=4.312e-12
+ PD=9.86e-06 PS=9.8e-07
mX57/X2/M0 N_X57/X2/8_X57/X2/M0_d N_STATE0_X57/X2/M0_g N_VSS_X57/X2/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=1.86e-12 PD=4.06e-06
+ PS=4.24e-06
mX57/X2/M1 N_X57/X2/10_X57/X2/M1_d N_X57/X2/8_X57/X2/M1_g N_VSS_X57/X2/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=7.95e-13 AS=1.5e-12 PD=5.3e-07
+ PS=4e-06
mX57/X2/M2 N_X57/X2/7_X57/X2/M2_d N_23_X57/X2/M2_g N_X57/X2/10_X57/X2/M2_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=7.95e-13 PD=4.06e-06
+ PS=5.3e-07
mX57/X2/M3 N_X57/X2/11_X57/X2/M3_d N_STATE0_X57/X2/M3_g N_VSS_X57/X2/M3_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=8.55e-13 AS=1.5e-12 PD=5.7e-07
+ PS=4e-06
mX57/X2/M4 N_X57/X2/9_X57/X2/M4_d N_INIT1_X57/X2/M4_g N_X57/X2/11_X57/X2/M4_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=8.55e-13 PD=4.08e-06
+ PS=5.7e-07
mX57/X2/M5 N_X57/X2/12_X57/X2/M5_d N_X57/X2/9_X57/X2/M5_g N_VSS_X57/X2/M5_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.86e-12 PD=9.8e-07
+ PS=4.24e-06
mX57/X2/M6 N_X57/11_X57/X2/M6_d N_X57/X2/7_X57/X2/M6_g N_X57/X2/12_X57/X2/M6_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=1.47e-12 PD=4.08e-06
+ PS=9.8e-07
mX57/X2/M7 N_X57/X2/8_X57/X2/M7_d N_STATE0_X57/X2/M7_g N_VDD_X57/X2/M7_s
+ N_VDD_X57/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=5.456e-12
+ PD=9.86e-06 PS=1.004e-05
mX57/X2/M8 N_X57/X2/7_X57/X2/M8_d N_X57/X2/8_X57/X2/M8_g N_VDD_X57/X2/M8_s
+ N_VDD_X57/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.332e-12 AS=4.4e-12 PD=5.3e-07
+ PS=9.8e-06
mX57/X2/M9 N_VDD_X57/X2/M9_d N_23_X57/X2/M9_g N_X57/X2/7_X57/X2/M9_s
+ N_VDD_X57/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=2.332e-12
+ PD=9.86e-06 PS=5.3e-07
mX57/X2/M10 N_X57/X2/9_X57/X2/M10_d N_STATE0_X57/X2/M10_g N_VDD_X57/X2/M10_s
+ N_VDD_X57/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.508e-12 AS=4.4e-12 PD=5.7e-07
+ PS=9.8e-06
mX57/X2/M11 N_VDD_X57/X2/M11_d N_INIT1_X57/X2/M11_g N_X57/X2/9_X57/X2/M11_s
+ N_VDD_X57/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=5.192e-12 AS=2.508e-12
+ PD=9.98e-06 PS=5.7e-07
mX57/X2/M12 N_X57/11_X57/X2/M12_d N_X57/X2/9_X57/X2/M12_g N_VDD_X57/X2/M12_s
+ N_VDD_X57/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.312e-12 AS=5.016e-12
+ PD=9.8e-07 PS=9.94e-06
mX57/X2/M13 N_VDD_X57/X2/M13_d N_X57/X2/7_X57/X2/M13_g N_X57/11_X57/X2/M13_s
+ N_VDD_X57/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=4.312e-12
+ PD=9.86e-06 PS=9.8e-07
mX58/X0/M0 N_X58/X0/8_X58/X0/M0_d N_STATE0_X58/X0/M0_g N_VSS_X58/X0/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=1.86e-12 PD=4.06e-06
+ PS=4.24e-06
mX58/X0/M1 N_X58/X0/10_X58/X0/M1_d N_X58/X0/8_X58/X0/M1_g N_VSS_X58/X0/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=7.95e-13 AS=1.5e-12 PD=5.3e-07
+ PS=4e-06
mX58/X0/M2 N_X58/X0/7_X58/X0/M2_d N_VSS_X58/X0/M2_g N_X58/X0/10_X58/X0/M2_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=7.95e-13 PD=4.06e-06
+ PS=5.3e-07
mX58/X0/M3 N_X58/X0/11_X58/X0/M3_d N_STATE0_X58/X0/M3_g N_VSS_X58/X0/M3_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=8.55e-13 AS=1.5e-12 PD=5.7e-07
+ PS=4e-06
mX58/X0/M4 N_X58/X0/9_X58/X0/M4_d N_VSS_X58/X0/M4_g N_X58/X0/11_X58/X0/M4_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=8.55e-13 PD=4.08e-06
+ PS=5.7e-07
mX58/X0/M5 N_X58/X0/12_X58/X0/M5_d N_X58/X0/9_X58/X0/M5_g N_VSS_X58/X0/M5_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.86e-12 PD=9.8e-07
+ PS=4.24e-06
mX58/X0/M6 N_X58/10_X58/X0/M6_d N_X58/X0/7_X58/X0/M6_g N_X58/X0/12_X58/X0/M6_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=1.47e-12 PD=4.08e-06
+ PS=9.8e-07
mX58/X0/M7 N_X58/X0/8_X58/X0/M7_d N_STATE0_X58/X0/M7_g N_VDD_X58/X0/M7_s
+ N_VDD_X58/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=5.456e-12
+ PD=9.86e-06 PS=1.004e-05
mX58/X0/M8 N_X58/X0/7_X58/X0/M8_d N_X58/X0/8_X58/X0/M8_g N_VDD_X58/X0/M8_s
+ N_VDD_X58/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.332e-12 AS=4.4e-12 PD=5.3e-07
+ PS=9.8e-06
mX58/X0/M9 N_VDD_X58/X0/M9_d N_VSS_X58/X0/M9_g N_X58/X0/7_X58/X0/M9_s
+ N_VDD_X58/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=2.332e-12
+ PD=9.86e-06 PS=5.3e-07
mX58/X0/M10 N_X58/X0/9_X58/X0/M10_d N_STATE0_X58/X0/M10_g N_VDD_X58/X0/M10_s
+ N_VDD_X58/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.508e-12 AS=4.4e-12 PD=5.7e-07
+ PS=9.8e-06
mX58/X0/M11 N_VDD_X58/X0/M11_d N_VSS_X58/X0/M11_g N_X58/X0/9_X58/X0/M11_s
+ N_VDD_X58/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=5.192e-12 AS=2.508e-12
+ PD=9.98e-06 PS=5.7e-07
mX58/X0/M12 N_X58/10_X58/X0/M12_d N_X58/X0/9_X58/X0/M12_g N_VDD_X58/X0/M12_s
+ N_VDD_X58/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.312e-12 AS=5.016e-12
+ PD=9.8e-07 PS=9.94e-06
mX58/X0/M13 N_VDD_X58/X0/M13_d N_X58/X0/7_X58/X0/M13_g N_X58/10_X58/X0/M13_s
+ N_VDD_X58/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=4.312e-12
+ PD=9.86e-06 PS=9.8e-07
mX58/X1/M0 N_X58/X1/8_X58/X1/M0_d N_STATE1_X58/X1/M0_g N_VSS_X58/X1/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=1.86e-12 PD=4.06e-06
+ PS=4.24e-06
mX58/X1/M1 N_X58/X1/10_X58/X1/M1_d N_X58/X1/8_X58/X1/M1_g N_VSS_X58/X1/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=7.95e-13 AS=1.5e-12 PD=5.3e-07
+ PS=4e-06
mX58/X1/M2 N_X58/X1/7_X58/X1/M2_d N_X58/10_X58/X1/M2_g N_X58/X1/10_X58/X1/M2_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=7.95e-13 PD=4.06e-06
+ PS=5.3e-07
mX58/X1/M3 N_X58/X1/11_X58/X1/M3_d N_STATE1_X58/X1/M3_g N_VSS_X58/X1/M3_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=8.55e-13 AS=1.5e-12 PD=5.7e-07
+ PS=4e-06
mX58/X1/M4 N_X58/X1/9_X58/X1/M4_d N_X58/11_X58/X1/M4_g N_X58/X1/11_X58/X1/M4_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=8.55e-13 PD=4.08e-06
+ PS=5.7e-07
mX58/X1/M5 N_X58/X1/12_X58/X1/M5_d N_X58/X1/9_X58/X1/M5_g N_VSS_X58/X1/M5_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.86e-12 PD=9.8e-07
+ PS=4.24e-06
mX58/X1/M6 N_MO3_X58/X1/M6_d N_X58/X1/7_X58/X1/M6_g N_X58/X1/12_X58/X1/M6_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=1.47e-12 PD=4.08e-06
+ PS=9.8e-07
mX58/X1/M7 N_X58/X1/8_X58/X1/M7_d N_STATE1_X58/X1/M7_g N_VDD_X58/X1/M7_s
+ N_VDD_X58/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=5.456e-12
+ PD=9.86e-06 PS=1.004e-05
mX58/X1/M8 N_X58/X1/7_X58/X1/M8_d N_X58/X1/8_X58/X1/M8_g N_VDD_X58/X1/M8_s
+ N_VDD_X58/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.332e-12 AS=4.4e-12 PD=5.3e-07
+ PS=9.8e-06
mX58/X1/M9 N_VDD_X58/X1/M9_d N_X58/10_X58/X1/M9_g N_X58/X1/7_X58/X1/M9_s
+ N_VDD_X58/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=2.332e-12
+ PD=9.86e-06 PS=5.3e-07
mX58/X1/M10 N_X58/X1/9_X58/X1/M10_d N_STATE1_X58/X1/M10_g N_VDD_X58/X1/M10_s
+ N_VDD_X58/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.508e-12 AS=4.4e-12 PD=5.7e-07
+ PS=9.8e-06
mX58/X1/M11 N_VDD_X58/X1/M11_d N_X58/11_X58/X1/M11_g N_X58/X1/9_X58/X1/M11_s
+ N_VDD_X58/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=5.192e-12 AS=2.508e-12
+ PD=9.98e-06 PS=5.7e-07
mX58/X1/M12 N_MO3_X58/X1/M12_d N_X58/X1/9_X58/X1/M12_g N_VDD_X58/X1/M12_s
+ N_VDD_X58/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.312e-12 AS=5.016e-12
+ PD=9.8e-07 PS=9.94e-06
mX58/X1/M13 N_VDD_X58/X1/M13_d N_X58/X1/7_X58/X1/M13_g N_MO3_X58/X1/M13_s
+ N_VDD_X58/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=4.312e-12
+ PD=9.86e-06 PS=9.8e-07
mX58/X2/M0 N_X58/X2/8_X58/X2/M0_d N_STATE0_X58/X2/M0_g N_VSS_X58/X2/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=1.86e-12 PD=4.06e-06
+ PS=4.24e-06
mX58/X2/M1 N_X58/X2/10_X58/X2/M1_d N_X58/X2/8_X58/X2/M1_g N_VSS_X58/X2/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=7.95e-13 AS=1.5e-12 PD=5.3e-07
+ PS=4e-06
mX58/X2/M2 N_X58/X2/7_X58/X2/M2_d N_14_X58/X2/M2_g N_X58/X2/10_X58/X2/M2_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=7.95e-13 PD=4.06e-06
+ PS=5.3e-07
mX58/X2/M3 N_X58/X2/11_X58/X2/M3_d N_STATE0_X58/X2/M3_g N_VSS_X58/X2/M3_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=8.55e-13 AS=1.5e-12 PD=5.7e-07
+ PS=4e-06
mX58/X2/M4 N_X58/X2/9_X58/X2/M4_d N_INIT3_X58/X2/M4_g N_X58/X2/11_X58/X2/M4_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=8.55e-13 PD=4.08e-06
+ PS=5.7e-07
mX58/X2/M5 N_X58/X2/12_X58/X2/M5_d N_X58/X2/9_X58/X2/M5_g N_VSS_X58/X2/M5_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.86e-12 PD=9.8e-07
+ PS=4.24e-06
mX58/X2/M6 N_X58/11_X58/X2/M6_d N_X58/X2/7_X58/X2/M6_g N_X58/X2/12_X58/X2/M6_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=1.47e-12 PD=4.08e-06
+ PS=9.8e-07
mX58/X2/M7 N_X58/X2/8_X58/X2/M7_d N_STATE0_X58/X2/M7_g N_VDD_X58/X2/M7_s
+ N_VDD_X58/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=5.456e-12
+ PD=9.86e-06 PS=1.004e-05
mX58/X2/M8 N_X58/X2/7_X58/X2/M8_d N_X58/X2/8_X58/X2/M8_g N_VDD_X58/X2/M8_s
+ N_VDD_X58/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.332e-12 AS=4.4e-12 PD=5.3e-07
+ PS=9.8e-06
mX58/X2/M9 N_VDD_X58/X2/M9_d N_14_X58/X2/M9_g N_X58/X2/7_X58/X2/M9_s
+ N_VDD_X58/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=2.332e-12
+ PD=9.86e-06 PS=5.3e-07
mX58/X2/M10 N_X58/X2/9_X58/X2/M10_d N_STATE0_X58/X2/M10_g N_VDD_X58/X2/M10_s
+ N_VDD_X58/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.508e-12 AS=4.4e-12 PD=5.7e-07
+ PS=9.8e-06
mX58/X2/M11 N_VDD_X58/X2/M11_d N_INIT3_X58/X2/M11_g N_X58/X2/9_X58/X2/M11_s
+ N_VDD_X58/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=5.192e-12 AS=2.508e-12
+ PD=9.98e-06 PS=5.7e-07
mX58/X2/M12 N_X58/11_X58/X2/M12_d N_X58/X2/9_X58/X2/M12_g N_VDD_X58/X2/M12_s
+ N_VDD_X58/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.312e-12 AS=5.016e-12
+ PD=9.8e-07 PS=9.94e-06
mX58/X2/M13 N_VDD_X58/X2/M13_d N_X58/X2/7_X58/X2/M13_g N_X58/11_X58/X2/M13_s
+ N_VDD_X58/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=4.312e-12
+ PD=9.86e-06 PS=9.8e-07
mX59/X0/M0 N_X59/X0/8_X59/X0/M0_d N_STATE0_X59/X0/M0_g N_VSS_X59/X0/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=1.86e-12 PD=4.06e-06
+ PS=4.24e-06
mX59/X0/M1 N_X59/X0/10_X59/X0/M1_d N_X59/X0/8_X59/X0/M1_g N_VSS_X59/X0/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=7.95e-13 AS=1.5e-12 PD=5.3e-07
+ PS=4e-06
mX59/X0/M2 N_X59/X0/7_X59/X0/M2_d N_VSS_X59/X0/M2_g N_X59/X0/10_X59/X0/M2_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=7.95e-13 PD=4.06e-06
+ PS=5.3e-07
mX59/X0/M3 N_X59/X0/11_X59/X0/M3_d N_STATE0_X59/X0/M3_g N_VSS_X59/X0/M3_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=8.55e-13 AS=1.5e-12 PD=5.7e-07
+ PS=4e-06
mX59/X0/M4 N_X59/X0/9_X59/X0/M4_d N_VSS_X59/X0/M4_g N_X59/X0/11_X59/X0/M4_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=8.55e-13 PD=4.08e-06
+ PS=5.7e-07
mX59/X0/M5 N_X59/X0/12_X59/X0/M5_d N_X59/X0/9_X59/X0/M5_g N_VSS_X59/X0/M5_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.86e-12 PD=9.8e-07
+ PS=4.24e-06
mX59/X0/M6 N_X59/10_X59/X0/M6_d N_X59/X0/7_X59/X0/M6_g N_X59/X0/12_X59/X0/M6_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=1.47e-12 PD=4.08e-06
+ PS=9.8e-07
mX59/X0/M7 N_X59/X0/8_X59/X0/M7_d N_STATE0_X59/X0/M7_g N_VDD_X59/X0/M7_s
+ N_VDD_X59/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=5.456e-12
+ PD=9.86e-06 PS=1.004e-05
mX59/X0/M8 N_X59/X0/7_X59/X0/M8_d N_X59/X0/8_X59/X0/M8_g N_VDD_X59/X0/M8_s
+ N_VDD_X59/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.332e-12 AS=4.4e-12 PD=5.3e-07
+ PS=9.8e-06
mX59/X0/M9 N_VDD_X59/X0/M9_d N_VSS_X59/X0/M9_g N_X59/X0/7_X59/X0/M9_s
+ N_VDD_X59/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=2.332e-12
+ PD=9.86e-06 PS=5.3e-07
mX59/X0/M10 N_X59/X0/9_X59/X0/M10_d N_STATE0_X59/X0/M10_g N_VDD_X59/X0/M10_s
+ N_VDD_X59/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.508e-12 AS=4.4e-12 PD=5.7e-07
+ PS=9.8e-06
mX59/X0/M11 N_VDD_X59/X0/M11_d N_VSS_X59/X0/M11_g N_X59/X0/9_X59/X0/M11_s
+ N_VDD_X59/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=5.192e-12 AS=2.508e-12
+ PD=9.98e-06 PS=5.7e-07
mX59/X0/M12 N_X59/10_X59/X0/M12_d N_X59/X0/9_X59/X0/M12_g N_VDD_X59/X0/M12_s
+ N_VDD_X59/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.312e-12 AS=5.016e-12
+ PD=9.8e-07 PS=9.94e-06
mX59/X0/M13 N_VDD_X59/X0/M13_d N_X59/X0/7_X59/X0/M13_g N_X59/10_X59/X0/M13_s
+ N_VDD_X59/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=4.312e-12
+ PD=9.86e-06 PS=9.8e-07
mX59/X1/M0 N_X59/X1/8_X59/X1/M0_d N_STATE1_X59/X1/M0_g N_VSS_X59/X1/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=1.86e-12 PD=4.06e-06
+ PS=4.24e-06
mX59/X1/M1 N_X59/X1/10_X59/X1/M1_d N_X59/X1/8_X59/X1/M1_g N_VSS_X59/X1/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=7.95e-13 AS=1.5e-12 PD=5.3e-07
+ PS=4e-06
mX59/X1/M2 N_X59/X1/7_X59/X1/M2_d N_X59/10_X59/X1/M2_g N_X59/X1/10_X59/X1/M2_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=7.95e-13 PD=4.06e-06
+ PS=5.3e-07
mX59/X1/M3 N_X59/X1/11_X59/X1/M3_d N_STATE1_X59/X1/M3_g N_VSS_X59/X1/M3_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=8.55e-13 AS=1.5e-12 PD=5.7e-07
+ PS=4e-06
mX59/X1/M4 N_X59/X1/9_X59/X1/M4_d N_X59/11_X59/X1/M4_g N_X59/X1/11_X59/X1/M4_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=8.55e-13 PD=4.08e-06
+ PS=5.7e-07
mX59/X1/M5 N_X59/X1/12_X59/X1/M5_d N_X59/X1/9_X59/X1/M5_g N_VSS_X59/X1/M5_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.86e-12 PD=9.8e-07
+ PS=4.24e-06
mX59/X1/M6 N_MO0_X59/X1/M6_d N_X59/X1/7_X59/X1/M6_g N_X59/X1/12_X59/X1/M6_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=1.47e-12 PD=4.08e-06
+ PS=9.8e-07
mX59/X1/M7 N_X59/X1/8_X59/X1/M7_d N_STATE1_X59/X1/M7_g N_VDD_X59/X1/M7_s
+ N_VDD_X59/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=5.456e-12
+ PD=9.86e-06 PS=1.004e-05
mX59/X1/M8 N_X59/X1/7_X59/X1/M8_d N_X59/X1/8_X59/X1/M8_g N_VDD_X59/X1/M8_s
+ N_VDD_X59/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.332e-12 AS=4.4e-12 PD=5.3e-07
+ PS=9.8e-06
mX59/X1/M9 N_VDD_X59/X1/M9_d N_X59/10_X59/X1/M9_g N_X59/X1/7_X59/X1/M9_s
+ N_VDD_X59/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=2.332e-12
+ PD=9.86e-06 PS=5.3e-07
mX59/X1/M10 N_X59/X1/9_X59/X1/M10_d N_STATE1_X59/X1/M10_g N_VDD_X59/X1/M10_s
+ N_VDD_X59/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.508e-12 AS=4.4e-12 PD=5.7e-07
+ PS=9.8e-06
mX59/X1/M11 N_VDD_X59/X1/M11_d N_X59/11_X59/X1/M11_g N_X59/X1/9_X59/X1/M11_s
+ N_VDD_X59/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=5.192e-12 AS=2.508e-12
+ PD=9.98e-06 PS=5.7e-07
mX59/X1/M12 N_MO0_X59/X1/M12_d N_X59/X1/9_X59/X1/M12_g N_VDD_X59/X1/M12_s
+ N_VDD_X59/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.312e-12 AS=5.016e-12
+ PD=9.8e-07 PS=9.94e-06
mX59/X1/M13 N_VDD_X59/X1/M13_d N_X59/X1/7_X59/X1/M13_g N_MO0_X59/X1/M13_s
+ N_VDD_X59/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=4.312e-12
+ PD=9.86e-06 PS=9.8e-07
mX59/X2/M0 N_X59/X2/8_X59/X2/M0_d N_STATE0_X59/X2/M0_g N_VSS_X59/X2/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=1.86e-12 PD=4.06e-06
+ PS=4.24e-06
mX59/X2/M1 N_X59/X2/10_X59/X2/M1_d N_X59/X2/8_X59/X2/M1_g N_VSS_X59/X2/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=7.95e-13 AS=1.5e-12 PD=5.3e-07
+ PS=4e-06
mX59/X2/M2 N_X59/X2/7_X59/X2/M2_d N_7_X59/X2/M2_g N_X59/X2/10_X59/X2/M2_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=7.95e-13 PD=4.06e-06
+ PS=5.3e-07
mX59/X2/M3 N_X59/X2/11_X59/X2/M3_d N_STATE0_X59/X2/M3_g N_VSS_X59/X2/M3_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=8.55e-13 AS=1.5e-12 PD=5.7e-07
+ PS=4e-06
mX59/X2/M4 N_X59/X2/9_X59/X2/M4_d N_INIT0_X59/X2/M4_g N_X59/X2/11_X59/X2/M4_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=8.55e-13 PD=4.08e-06
+ PS=5.7e-07
mX59/X2/M5 N_X59/X2/12_X59/X2/M5_d N_X59/X2/9_X59/X2/M5_g N_VSS_X59/X2/M5_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.86e-12 PD=9.8e-07
+ PS=4.24e-06
mX59/X2/M6 N_X59/11_X59/X2/M6_d N_X59/X2/7_X59/X2/M6_g N_X59/X2/12_X59/X2/M6_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=1.47e-12 PD=4.08e-06
+ PS=9.8e-07
mX59/X2/M7 N_X59/X2/8_X59/X2/M7_d N_STATE0_X59/X2/M7_g N_VDD_X59/X2/M7_s
+ N_VDD_X59/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=5.456e-12
+ PD=9.86e-06 PS=1.004e-05
mX59/X2/M8 N_X59/X2/7_X59/X2/M8_d N_X59/X2/8_X59/X2/M8_g N_VDD_X59/X2/M8_s
+ N_VDD_X59/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.332e-12 AS=4.4e-12 PD=5.3e-07
+ PS=9.8e-06
mX59/X2/M9 N_VDD_X59/X2/M9_d N_7_X59/X2/M9_g N_X59/X2/7_X59/X2/M9_s
+ N_VDD_X59/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=2.332e-12
+ PD=9.86e-06 PS=5.3e-07
mX59/X2/M10 N_X59/X2/9_X59/X2/M10_d N_STATE0_X59/X2/M10_g N_VDD_X59/X2/M10_s
+ N_VDD_X59/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.508e-12 AS=4.4e-12 PD=5.7e-07
+ PS=9.8e-06
mX59/X2/M11 N_VDD_X59/X2/M11_d N_INIT0_X59/X2/M11_g N_X59/X2/9_X59/X2/M11_s
+ N_VDD_X59/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=5.192e-12 AS=2.508e-12
+ PD=9.98e-06 PS=5.7e-07
mX59/X2/M12 N_X59/11_X59/X2/M12_d N_X59/X2/9_X59/X2/M12_g N_VDD_X59/X2/M12_s
+ N_VDD_X59/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.312e-12 AS=5.016e-12
+ PD=9.8e-07 PS=9.94e-06
mX59/X2/M13 N_VDD_X59/X2/M13_d N_X59/X2/7_X59/X2/M13_g N_X59/11_X59/X2/M13_s
+ N_VDD_X59/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=4.312e-12
+ PD=9.86e-06 PS=9.8e-07
mX60/X0/M0 N_X60/X0/8_X60/X0/M0_d N_STATE0_X60/X0/M0_g N_VSS_X60/X0/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=1.86e-12 PD=4.06e-06
+ PS=4.24e-06
mX60/X0/M1 N_X60/X0/10_X60/X0/M1_d N_X60/X0/8_X60/X0/M1_g N_VSS_X60/X0/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=7.95e-13 AS=1.5e-12 PD=5.3e-07
+ PS=4e-06
mX60/X0/M2 N_X60/X0/7_X60/X0/M2_d N_VSS_X60/X0/M2_g N_X60/X0/10_X60/X0/M2_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=7.95e-13 PD=4.06e-06
+ PS=5.3e-07
mX60/X0/M3 N_X60/X0/11_X60/X0/M3_d N_STATE0_X60/X0/M3_g N_VSS_X60/X0/M3_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=8.55e-13 AS=1.5e-12 PD=5.7e-07
+ PS=4e-06
mX60/X0/M4 N_X60/X0/9_X60/X0/M4_d N_VSS_X60/X0/M4_g N_X60/X0/11_X60/X0/M4_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=8.55e-13 PD=4.08e-06
+ PS=5.7e-07
mX60/X0/M5 N_X60/X0/12_X60/X0/M5_d N_X60/X0/9_X60/X0/M5_g N_VSS_X60/X0/M5_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.86e-12 PD=9.8e-07
+ PS=4.24e-06
mX60/X0/M6 N_X60/10_X60/X0/M6_d N_X60/X0/7_X60/X0/M6_g N_X60/X0/12_X60/X0/M6_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=1.47e-12 PD=4.08e-06
+ PS=9.8e-07
mX60/X0/M7 N_X60/X0/8_X60/X0/M7_d N_STATE0_X60/X0/M7_g N_VDD_X60/X0/M7_s
+ N_VDD_X60/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=5.456e-12
+ PD=9.86e-06 PS=1.004e-05
mX60/X0/M8 N_X60/X0/7_X60/X0/M8_d N_X60/X0/8_X60/X0/M8_g N_VDD_X60/X0/M8_s
+ N_VDD_X60/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.332e-12 AS=4.4e-12 PD=5.3e-07
+ PS=9.8e-06
mX60/X0/M9 N_VDD_X60/X0/M9_d N_VSS_X60/X0/M9_g N_X60/X0/7_X60/X0/M9_s
+ N_VDD_X60/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=2.332e-12
+ PD=9.86e-06 PS=5.3e-07
mX60/X0/M10 N_X60/X0/9_X60/X0/M10_d N_STATE0_X60/X0/M10_g N_VDD_X60/X0/M10_s
+ N_VDD_X60/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.508e-12 AS=4.4e-12 PD=5.7e-07
+ PS=9.8e-06
mX60/X0/M11 N_VDD_X60/X0/M11_d N_VSS_X60/X0/M11_g N_X60/X0/9_X60/X0/M11_s
+ N_VDD_X60/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=5.192e-12 AS=2.508e-12
+ PD=9.98e-06 PS=5.7e-07
mX60/X0/M12 N_X60/10_X60/X0/M12_d N_X60/X0/9_X60/X0/M12_g N_VDD_X60/X0/M12_s
+ N_VDD_X60/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.312e-12 AS=5.016e-12
+ PD=9.8e-07 PS=9.94e-06
mX60/X0/M13 N_VDD_X60/X0/M13_d N_X60/X0/7_X60/X0/M13_g N_X60/10_X60/X0/M13_s
+ N_VDD_X60/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=4.312e-12
+ PD=9.86e-06 PS=9.8e-07
mX60/X1/M0 N_X60/X1/8_X60/X1/M0_d N_STATE1_X60/X1/M0_g N_VSS_X60/X1/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=1.86e-12 PD=4.06e-06
+ PS=4.24e-06
mX60/X1/M1 N_X60/X1/10_X60/X1/M1_d N_X60/X1/8_X60/X1/M1_g N_VSS_X60/X1/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=7.95e-13 AS=1.5e-12 PD=5.3e-07
+ PS=4e-06
mX60/X1/M2 N_X60/X1/7_X60/X1/M2_d N_X60/10_X60/X1/M2_g N_X60/X1/10_X60/X1/M2_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=7.95e-13 PD=4.06e-06
+ PS=5.3e-07
mX60/X1/M3 N_X60/X1/11_X60/X1/M3_d N_STATE1_X60/X1/M3_g N_VSS_X60/X1/M3_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=8.55e-13 AS=1.5e-12 PD=5.7e-07
+ PS=4e-06
mX60/X1/M4 N_X60/X1/9_X60/X1/M4_d N_X60/11_X60/X1/M4_g N_X60/X1/11_X60/X1/M4_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=8.55e-13 PD=4.08e-06
+ PS=5.7e-07
mX60/X1/M5 N_X60/X1/12_X60/X1/M5_d N_X60/X1/9_X60/X1/M5_g N_VSS_X60/X1/M5_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.86e-12 PD=9.8e-07
+ PS=4.24e-06
mX60/X1/M6 N_MO2_X60/X1/M6_d N_X60/X1/7_X60/X1/M6_g N_X60/X1/12_X60/X1/M6_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=1.47e-12 PD=4.08e-06
+ PS=9.8e-07
mX60/X1/M7 N_X60/X1/8_X60/X1/M7_d N_STATE1_X60/X1/M7_g N_VDD_X60/X1/M7_s
+ N_VDD_X60/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=5.456e-12
+ PD=9.86e-06 PS=1.004e-05
mX60/X1/M8 N_X60/X1/7_X60/X1/M8_d N_X60/X1/8_X60/X1/M8_g N_VDD_X60/X1/M8_s
+ N_VDD_X60/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.332e-12 AS=4.4e-12 PD=5.3e-07
+ PS=9.8e-06
mX60/X1/M9 N_VDD_X60/X1/M9_d N_X60/10_X60/X1/M9_g N_X60/X1/7_X60/X1/M9_s
+ N_VDD_X60/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=2.332e-12
+ PD=9.86e-06 PS=5.3e-07
mX60/X1/M10 N_X60/X1/9_X60/X1/M10_d N_STATE1_X60/X1/M10_g N_VDD_X60/X1/M10_s
+ N_VDD_X60/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.508e-12 AS=4.4e-12 PD=5.7e-07
+ PS=9.8e-06
mX60/X1/M11 N_VDD_X60/X1/M11_d N_X60/11_X60/X1/M11_g N_X60/X1/9_X60/X1/M11_s
+ N_VDD_X60/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=5.192e-12 AS=2.508e-12
+ PD=9.98e-06 PS=5.7e-07
mX60/X1/M12 N_MO2_X60/X1/M12_d N_X60/X1/9_X60/X1/M12_g N_VDD_X60/X1/M12_s
+ N_VDD_X60/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.312e-12 AS=5.016e-12
+ PD=9.8e-07 PS=9.94e-06
mX60/X1/M13 N_VDD_X60/X1/M13_d N_X60/X1/7_X60/X1/M13_g N_MO2_X60/X1/M13_s
+ N_VDD_X60/X1/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=4.312e-12
+ PD=9.86e-06 PS=9.8e-07
mX60/X2/M0 N_X60/X2/8_X60/X2/M0_d N_STATE0_X60/X2/M0_g N_VSS_X60/X2/M0_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=1.86e-12 PD=4.06e-06
+ PS=4.24e-06
mX60/X2/M1 N_X60/X2/10_X60/X2/M1_d N_X60/X2/8_X60/X2/M1_g N_VSS_X60/X2/M1_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=7.95e-13 AS=1.5e-12 PD=5.3e-07
+ PS=4e-06
mX60/X2/M2 N_X60/X2/7_X60/X2/M2_d N_20_X60/X2/M2_g N_X60/X2/10_X60/X2/M2_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.59e-12 AS=7.95e-13 PD=4.06e-06
+ PS=5.3e-07
mX60/X2/M3 N_X60/X2/11_X60/X2/M3_d N_STATE0_X60/X2/M3_g N_VSS_X60/X2/M3_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=8.55e-13 AS=1.5e-12 PD=5.7e-07
+ PS=4e-06
mX60/X2/M4 N_X60/X2/9_X60/X2/M4_d N_INIT2_X60/X2/M4_g N_X60/X2/11_X60/X2/M4_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=8.55e-13 PD=4.08e-06
+ PS=5.7e-07
mX60/X2/M5 N_X60/X2/12_X60/X2/M5_d N_X60/X2/9_X60/X2/M5_g N_VSS_X60/X2/M5_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.86e-12 PD=9.8e-07
+ PS=4.24e-06
mX60/X2/M6 N_X60/11_X60/X2/M6_d N_X60/X2/7_X60/X2/M6_g N_X60/X2/12_X60/X2/M6_s
+ N_VSS_X24/M0_b N_18 L=1.8e-07 W=3e-06 AD=1.62e-12 AS=1.47e-12 PD=4.08e-06
+ PS=9.8e-07
mX60/X2/M7 N_X60/X2/8_X60/X2/M7_d N_STATE0_X60/X2/M7_g N_VDD_X60/X2/M7_s
+ N_VDD_X60/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=5.456e-12
+ PD=9.86e-06 PS=1.004e-05
mX60/X2/M8 N_X60/X2/7_X60/X2/M8_d N_X60/X2/8_X60/X2/M8_g N_VDD_X60/X2/M8_s
+ N_VDD_X60/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.332e-12 AS=4.4e-12 PD=5.3e-07
+ PS=9.8e-06
mX60/X2/M9 N_VDD_X60/X2/M9_d N_20_X60/X2/M9_g N_X60/X2/7_X60/X2/M9_s
+ N_VDD_X60/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=2.332e-12
+ PD=9.86e-06 PS=5.3e-07
mX60/X2/M10 N_X60/X2/9_X60/X2/M10_d N_STATE0_X60/X2/M10_g N_VDD_X60/X2/M10_s
+ N_VDD_X60/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=2.508e-12 AS=4.4e-12 PD=5.7e-07
+ PS=9.8e-06
mX60/X2/M11 N_VDD_X60/X2/M11_d N_INIT2_X60/X2/M11_g N_X60/X2/9_X60/X2/M11_s
+ N_VDD_X60/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=5.192e-12 AS=2.508e-12
+ PD=9.98e-06 PS=5.7e-07
mX60/X2/M12 N_X60/11_X60/X2/M12_d N_X60/X2/9_X60/X2/M12_g N_VDD_X60/X2/M12_s
+ N_VDD_X60/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.312e-12 AS=5.016e-12
+ PD=9.8e-07 PS=9.94e-06
mX60/X2/M13 N_VDD_X60/X2/M13_d N_X60/X2/7_X60/X2/M13_g N_X60/11_X60/X2/M13_s
+ N_VDD_X60/X0/M7_b P_18 L=1.8e-07 W=8.8e-06 AD=4.664e-12 AS=4.312e-12
+ PD=9.86e-06 PS=9.8e-07
*
.include "Coin_bank.pex.sp.COIN_BANK.pxi"
*
.ends
*
*
